`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Dr.EDWIN DHAS D
// 
// Create Date: 02.10.2024 13:11:01
// Design Name: 
// Module Name: adding_8
// Project Name: CNN-based digit classification 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module main_program #(parameter w1=10, parameter w2=21, parameter w3=9, parameter w4=18, parameter w5=10, parameter w6=21, parameter w7=18, parameter w8=24, parameter w9=9, parameter w10=10, parameter w11=21, parameter w12=27, parameter w13=18, parameter w14=9, parameter w15=64)(
input clk,
input rst,
input signed [8:0] inp,
output signed [w2-1: 0] oup1, oup2, oup3, oup4, oup5, oup6, oup7, oup8,
output signed [w8-1:0] add1, add2, add3, add4,add5,add6,add7, add8,add9, add10, add11, add12,add13,add14,add15, add16,
output signed [w12-1:0] ad1,ad2,ad3,ad4,ad5,ad6,ad7,ad8,ad9,ad10,ad11,ad12,ad13,ad14,ad15,ad16,ad17,ad18,ad19,ad20,ad21,ad22,ad23,ad24,ad25,ad26,ad27,ad28,ad29,ad30,ad31,ad32,
output En1,En9, En137,enf,
output clk1,clk3,
output [3:0] max_index
    );


wire [w15-1:0] op1,op2, op3, op4, op5,op6,op7, op8, op9, op10;
wire [w15-1:0] oc1,oc2, oc3, oc4, oc5,oc6,oc7, oc8, oc9, oc10;
//wire enf;
//wire max_index;
wire En2, En3, En4, En5, En6, En7, En8;
//wire signed [w2-1: 0] oup1, oup2, oup3, oup4, oup5, oup6, oup7, oup8;
wire signed [w3-1:0] ou1,ou2,ou3,ou4,ou5,ou6,ou7,ou8;
wire signed [w3-1:0] oua1,oua2,oua3,oua4,oua5,oua6,oua7,oua8;
wire signed [w3-1:0] ouy1,ouy2,ouy3,ouy4,ouy5,ouy6,ouy7,ouy8;
reg signed [w3-1:0] ouz1,ouz2,ouz3,ouz4,ouz5,ouz6,ouz7,ouz8;
reg signed [w3-1:0] oux1,oux2,oux3,oux4,oux5,oux6,oux7,oux8;
wire E10,E11,E12,E13,E14, E15, E16, E17;
wire signed [w3-1:0] oub1,oub2,oub3,oub4,oub5,oub6,oub7,oub8;
reg Ea=1'b0;
reg Eb=1'b0;
wire signed [w6-1:0] oup9, oup10, oup11, oup12, oup13, oup14, oup15, oup16, oup17, oup18, oup19, oup20, oup21, oup22, oup23, oup24, oup25, oup26, oup27, oup28, oup29, oup30, oup31, oup32, oup33, oup34, oup35, oup36, oup37, oup38, oup39, oup40, oup41, oup42, oup43, oup44, oup45, oup46, oup47, oup48, oup49, oup50, oup51, oup52, oup53, oup54, oup55, oup56, oup57, oup58, oup59, oup60, oup61, oup62, oup63, oup64, oup65, oup66, oup67, oup68, oup69, oup70, oup71, oup72, oup73, oup74, oup75, oup76, oup77, oup78, oup79, oup80, oup81, oup82, oup83, oup84, oup85, oup86, oup87, oup88, oup89, oup90, oup91, oup92, oup93, oup94, oup95, oup96, oup97, oup98, oup99, oup100, oup101, oup102, oup103, oup104, oup105, oup106, oup107, oup108, oup109, oup110, oup111, oup112, oup113, oup114, oup115, oup116, oup117, oup118, oup119, oup120, oup121, oup122, oup123, oup124, oup125, oup126, oup127, oup128, oup129, oup130, oup131, oup132, oup133, oup134, oup135, oup136;
//wire signed [w8-1:0] add1, add2, add3, add4,add5,add6,add7, add8,add9, add10, add11, add12,add13,add14,add15, add16;
reg rst1=1'b1;
reg rst3=1'b1;
reg rst4=1'b1;
wire  En10,  En11,  En12,  En13,  En14,  En15,  En16,  En17,  En18,  En19,  En20,  En21,  En22,  En23,  En24,  En25,  En26,  En27,  En28,  En29,  En30,  En31,  En32,  En33,  En34,  En35,  En36,  En37,  En38,  En39,  En40,  En41,  En42,  En43,  En44,  En45,  En46,  En47,  En48,  En49,  En50,  En51,  En52,  En53,  En54,  En55,  En56,  En57,  En58,  En59,  En60,  En61,  En62,  En63,  En64,  En65,  En66,  En67,  En68,  En69,  En70,  En71,  En72,  En73,  En74,  En75,  En76,  En77,  En78,  En79,  En80,  En81,  En82,  En83,  En84,  En85,  En86,  En87,  En88,  En89,  En90,  En91,  En92,  En93,  En94,  En95,  En96,  En97,  En98,  En99,  En100,  En101,  En102,  En103,  En104,  En105,  En106,  En107,  En108,  En109,  En110,  En111,  En112,  En113,  En114,  En115,  En116,  En117,  En118,  En119,  En120,  En121,  En122,  En123,  En124,  En125,  En126,  En127,  En128,  En129,  En130,  En131,  En132,  En133,  En134,  En135,  En136;
//wire clk1;
//wire clk3;
wire [w9-1:0] bn_ou1, bn_ou2,bn_ou3, bn_ou4,bn_ou5, bn_ou6,bn_ou7,bn_ou8,bn_ou9, bn_ou10,bn_ou11, bn_ou12,bn_ou13, bn_ou14,bn_ou15,bn_ou16;
wire [w9-1:0] ro1,ro2,ro3,ro4,ro5,ro6,ro7,ro8,ro9,ro10,ro11,ro12,ro13,ro14,ro15,ro16;
wire enab1,enab2,enab3,enab4,enab5,enab6,enab7,enab8,enab9,enab10,enab11,enab12,enab13,enab14,enab15,enab16;
wire [w9-1:0] mp_ou1,mp_ou2,mp_ou3,mp_ou4,mp_ou5,mp_ou6,mp_ou7,mp_ou8,mp_ou9,mp_ou10,mp_ou11,mp_ou12,mp_ou13,mp_ou14,mp_ou15,mp_ou16;
reg [w9-1:0] roa1,roa2,roa3,roa4,roa5,roa6,roa7,roa8,roa9,roa10,roa11,roa12,roa13,roa14,roa15,roa16;
wire  En138,  En139,  En140,  En141,  En142,  En143,  En144,  En145,  En146,  En147,  En148,  En149,  En150,  En151,  En152,  En153,  En154,  En155,  En156,  En157,  En158,  En159,  En160,  En161,  En162,  En163,  En164,  En165,  En166,  En167,  En168,  En169,  En170,  En171,  En172,  En173,  En174,  En175,  En176,  En177,  En178,  En179,  En180,  En181,  En182,  En183,  En184,  En185,  En186,  En187,  En188,  En189,  En190,  En191,  En192,  En193,  En194,  En195,  En196,  En197,  En198,  En199,  En200,  En201,  En202,  En203,  En204,  En205,  En206,  En207,  En208,  En209,  En210,  En211,  En212,  En213,  En214,  En215,  En216,  En217,  En218,  En219,  En220,  En221,  En222,  En223,  En224,  En225,  En226,  En227,  En228,  En229,  En230,  En231,  En232,  En233,  En234,  En235,  En236,  En237,  En238,  En239,  En240,  En241,  En242,  En243,  En244,  En245,  En246,  En247,  En248,  En249,  En250,  En251,  En252,  En253,  En254,  En255,  En256,  En257,  En258,  En259,  En260,  En261,  En262,  En263,  En264,  En265,  En266,  En267,  En268,  En269,  En270,  En271,  En272,  En273,  En274,  En275,  En276,  En277,  En278,  En279,  En280,  En281,  En282,  En283,  En284,  En285,  En286,  En287,  En288,  En289,  En290,  En291,  En292,  En293,  En294,  En295,  En296,  En297,  En298,  En299,  En300,  En301,  En302,  En303,  En304,  En305,  En306,  En307,  En308,  En309,  En310,  En311,  En312,  En313,  En314,  En315,  En316,  En317,  En318,  En319,  En320,  En321,  En322,  En323,  En324,  En325,  En326,  En327,  En328,  En329,  En330,  En331,  En332,  En333,  En334,  En335,  En336,  En337,  En338,  En339,  En340,  En341,  En342,  En343,  En344,  En345,  En346,  En347,  En348,  En349,  En350,  En351,  En352,  En353,  En354,  En355,  En356,  En357,  En358,  En359,  En360,  En361,  En362,  En363,  En364,  En365,  En366,  En367,  En368,  En369,  En370,  En371,  En372,  En373,  En374,  En375,  En376,  En377,  En378,  En379,  En380,  En381,  En382,  En383,  En384,  En385,  En386,  En387,  En388,  En389,  En390,  En391,  En392,  En393,  En394,  En395,  En396,  En397,  En398,  En399,  En400,  En401,  En402,  En403,  En404,  En405,  En406,  En407,  En408,  En409,  En410,  En411,  En412,  En413,  En414,  En415,  En416,  En417,  En418,  En419,  En420,  En421,  En422,  En423,  En424,  En425,  En426,  En427,  En428,  En429,  En430,  En431,  En432,  En433,  En434,  En435,  En436,  En437,  En438,  En439,  En440,  En441,  En442,  En443,  En444,  En445,  En446,  En447,  En448,  En449,  En450,  En451,  En452,  En453,  En454,  En455,  En456,  En457,  En458,  En459,  En460,  En461,  En462,  En463,  En464,  En465,  En466,  En467,  En468,  En469,  En470,  En471,  En472,  En473,  En474,  En475,  En476,  En477,  En478,  En479,  En480,  En481,  En482,  En483,  En484,  En485,  En486,  En487,  En488,  En489,  En490,  En491,  En492,  En493,  En494,  En495,  En496,  En497,  En498,  En499,  En500,  En501,  En502,  En503,  En504,  En505,  En506,  En507,  En508,  En509,  En510,  En511,  En512,  En513,  En514,  En515,  En516,  En517,  En518,  En519,  En520,  En521,  En522,  En523,  En524,  En525,  En526,  En527,  En528,  En529,  En530,  En531,  En532,  En533,  En534,  En535,  En536,  En537,  En538,  En539,  En540,  En541,  En542,  En543,  En544,  En545,  En546,  En547,  En548,  En549,  En550,  En551,  En552,  En553,  En554,  En555,  En556,  En557,  En558,  En559,  En560,  En561,  En562,  En563,  En564,  En565,  En566,  En567,  En568,  En569,  En570,  En571,  En572,  En573,  En574,  En575,  En576,  En577,  En578,  En579,  En580,  En581,  En582,  En583,  En584,  En585,  En586,  En587,  En588,  En589,  En590,  En591,  En592,  En593,  En594,  En595,  En596,  En597,  En598,  En599,  En600,  En601,  En602,  En603,  En604,  En605,  En606,  En607,  En608,  En609,  En610,  En611,  En612,  En613,  En614,  En615,  En616,  En617,  En618,  En619,  En620,  En621,  En622,  En623,  En624,  En625,  En626,  En627,  En628,  En629,  En630,  En631,  En632,  En633,  En634,  En635,  En636,  En637,  En638,  En639,  En640,  En641,  En642,  En643,  En644,  En645,  En646,  En647,  En648;


wire [w14-1:0] bn_ou17,bn_ou18,bn_ou19,bn_ou20,bn_ou21,bn_ou22,bn_ou23,bn_ou24,bn_ou25,bn_ou26,bn_ou27,bn_ou28,bn_ou29,bn_ou30,bn_ou31,bn_ou32,bn_ou33,bn_ou34,bn_ou35,bn_ou36,bn_ou37,bn_ou38,bn_ou39,bn_ou40,bn_ou41,bn_ou42,bn_ou43,bn_ou44,bn_ou45,bn_ou46,bn_ou47,bn_ou48;
wire   [w14-1:0] ro17, ro18,ro19, ro20,ro21, ro22,ro23, ro24,ro25, ro26,ro27, ro28,ro29, ro30,ro31, ro32,ro33, ro34,ro35, ro36,ro37, ro38,ro39, ro40,ro41, ro42,ro43, ro44,ro45, ro46,ro47, ro48;

wire [w11-1:0] oud137, oud138, oud139, oud140, oud141, oud142, oud143, oud144, oud145, oud146, oud147, oud148, oud149, oud150, oud151, oud152, oud153, oud154, oud155, oud156, oud157, oud158, oud159, oud160, oud161, oud162, oud163, oud164, oud165, oud166, oud167, oud168, oud169, oud170, oud171, oud172, oud173, oud174, oud175, oud176, oud177, oud178, oud179, oud180, oud181, oud182, oud183, oud184, oud185, oud186, oud187, oud188, oud189, oud190, oud191, oud192, oud193, oud194, oud195, oud196, oud197, oud198, oud199, oud200, oud201, oud202, oud203, oud204, oud205, oud206, oud207, oud208, oud209, oud210, oud211, oud212, oud213, oud214, oud215, oud216, oud217, oud218, oud219, oud220, oud221, oud222, oud223, oud224, oud225, oud226, oud227, oud228, oud229, oud230, oud231, oud232, oud233, oud234, oud235, oud236, oud237, oud238, oud239, oud240, oud241, oud242, oud243, oud244, oud245, oud246, oud247, oud248, oud249, oud250, oud251, oud252, oud253, oud254, oud255, oud256, oud257, oud258, oud259, oud260, oud261, oud262, oud263, oud264, oud265, oud266, oud267, oud268, oud269, oud270, oud271, oud272, oud273, oud274, oud275, oud276, oud277, oud278, oud279, oud280, oud281, oud282, oud283, oud284, oud285, oud286, oud287, oud288, oud289, oud290, oud291, oud292, oud293, oud294, oud295, oud296, oud297, oud298, oud299, oud300, oud301, oud302, oud303, oud304, oud305, oud306, oud307, oud308, oud309, oud310, oud311, oud312, oud313, oud314, oud315, oud316, oud317, oud318, oud319, oud320, oud321, oud322, oud323, oud324, oud325, oud326, oud327, oud328, oud329, oud330, oud331, oud332, oud333, oud334, oud335, oud336, oud337, oud338, oud339, oud340, oud341, oud342, oud343, oud344, oud345, oud346, oud347, oud348, oud349, oud350, oud351, oud352, oud353, oud354, oud355, oud356, oud357, oud358, oud359, oud360, oud361, oud362, oud363, oud364, oud365, oud366, oud367, oud368, oud369, oud370, oud371, oud372, oud373, oud374, oud375, oud376, oud377, oud378, oud379, oud380, oud381, oud382, oud383, oud384, oud385, oud386, oud387, oud388, oud389, oud390, oud391, oud392, oud393, oud394, oud395, oud396, oud397, oud398, oud399, oud400, oud401, oud402, oud403, oud404, oud405, oud406, oud407, oud408, oud409, oud410, oud411, oud412, oud413, oud414, oud415, oud416, oud417, oud418, oud419, oud420, oud421, oud422, oud423, oud424, oud425, oud426, oud427, oud428, oud429, oud430, oud431, oud432, oud433, oud434, oud435, oud436, oud437, oud438, oud439, oud440, oud441, oud442, oud443, oud444, oud445, oud446, oud447, oud448, oud449, oud450, oud451, oud452, oud453, oud454, oud455, oud456, oud457, oud458, oud459, oud460, oud461, oud462, oud463, oud464, oud465, oud466, oud467, oud468, oud469, oud470, oud471, oud472, oud473, oud474, oud475, oud476, oud477, oud478, oud479, oud480, oud481, oud482, oud483, oud484, oud485, oud486, oud487, oud488, oud489, oud490, oud491, oud492, oud493, oud494, oud495, oud496, oud497, oud498, oud499, oud500, oud501, oud502, oud503, oud504, oud505, oud506, oud507, oud508, oud509, oud510, oud511, oud512, oud513, oud514, oud515, oud516, oud517, oud518, oud519, oud520, oud521, oud522, oud523, oud524, oud525, oud526, oud527, oud528, oud529, oud530, oud531, oud532, oud533, oud534, oud535, oud536, oud537, oud538, oud539, oud540, oud541, oud542, oud543, oud544, oud545, oud546, oud547, oud548, oud549, oud550, oud551, oud552, oud553, oud554, oud555, oud556, oud557, oud558, oud559, oud560, oud561, oud562, oud563, oud564, oud565, oud566, oud567, oud568, oud569, oud570, oud571, oud572, oud573, oud574, oud575, oud576, oud577, oud578, oud579, oud580, oud581, oud582, oud583, oud584, oud585, oud586, oud587, oud588, oud589, oud590, oud591, oud592, oud593, oud594, oud595, oud596, oud597, oud598, oud599, oud600, oud601, oud602, oud603, oud604, oud605, oud606, oud607, oud608, oud609, oud610, oud611, oud612, oud613, oud614, oud615, oud616, oud617, oud618, oud619, oud620, oud621, oud622, oud623, oud624, oud625, oud626, oud627, oud628, oud629, oud630, oud631, oud632, oud633, oud634, oud635, oud636, oud637, oud638, oud639, oud640, oud641, oud642, oud643, oud644, oud645, oud646, oud647, oud648;
//wire [w12-1:0] ad1,ad2,ad3,ad4,ad5,ad6,ad7,ad8,ad9,ad10,ad11,ad12,ad13,ad14,ad15,ad16,ad17,ad18,ad19,ad20,ad21,ad22,ad23,ad24,ad25,ad26,ad27,ad28,ad29,ad30,ad31,ad32;
reg [w9-1:0] ouf1,ouf2,ouf3, ouf4,ouf5,ouf6,ouf7, ouf8,ouf9,ouf10,ouf11, ouf12,ouf13,ouf14,ouf15, ouf16;
reg [w14-1:0] r17, r18,r19, r20,r21, r22,r23, r24,r25, r26,r27, r28,r29, r30,r31, r32,r33, r34,r35, r36,r37, r38,r39, r40,r41, r42,r43, r44,r45, r46,r47, r48;
wire f_en;
wire [w14-1:0] f_ou;
reg [w14-1:0] f_ou1;
reg rst5=1'b1;
//wire [3:0] max_index;

//assign ouv=f_ou;


//assign En=enf;
//assign clk_out=clk3;
reg signed [w1-1:0] ka1=125;	reg signed [w1-1:0] kb1=87;	reg signed [w1-1:0] kc1=-212;	reg signed [w1-1:0] kd1=211;	reg signed [w1-1:0] ke1=-170;	reg signed [w1-1:0] kf1=-77;	reg signed [w1-1:0] kg1=-9;	reg signed [w1-1:0] kh1=-175;	reg signed [w1-1:0] ki1=-167;
reg signed [w1-1:0] ka2=-73;	reg signed [w1-1:0] kb2=-30;	reg signed [w1-1:0] kc2=-26;	reg signed [w1-1:0] kd2=-153;	reg signed [w1-1:0] ke2=-314;	reg signed [w1-1:0] kf2=-214;	reg signed [w1-1:0] kg2=249;	reg signed [w1-1:0] kh2=305;	reg signed [w1-1:0] ki2=72;
reg signed [w1-1:0] ka3=279;	reg signed [w1-1:0] kb3=-177;	reg signed [w1-1:0] kc3=-24;	reg signed [w1-1:0] kd3=209;	reg signed [w1-1:0] ke3=-150;	reg signed [w1-1:0] kf3=201;	reg signed [w1-1:0] kg3=7;	reg signed [w1-1:0] kh3=35;	reg signed [w1-1:0] ki3=-314;
reg signed [w1-1:0] ka4=104;	reg signed [w1-1:0] kb4=30;	reg signed [w1-1:0] kc4=233;	reg signed [w1-1:0] kd4=-91;	reg signed [w1-1:0] ke4=300;	reg signed [w1-1:0] kf4=-313;	reg signed [w1-1:0] kg4=-98;	reg signed [w1-1:0] kh4=261;	reg signed [w1-1:0] ki4=-161;
reg signed [w1-1:0] ka5=320;	reg signed [w1-1:0] kb5=223;	reg signed [w1-1:0] kc5=-269;	reg signed [w1-1:0] kd5=-308;	reg signed [w1-1:0] ke5=-251;	reg signed [w1-1:0] kf5=-76;	reg signed [w1-1:0] kg5=33;	reg signed [w1-1:0] kh5=197;	reg signed [w1-1:0] ki5=-65;
reg signed [w1-1:0] ka6=330;	reg signed [w1-1:0] kb6=134;	reg signed [w1-1:0] kc6=-158;	reg signed [w1-1:0] kd6=120;	reg signed [w1-1:0] ke6=148;	reg signed [w1-1:0] kf6=120;	reg signed [w1-1:0] kg6=108;	reg signed [w1-1:0] kh6=199;	reg signed [w1-1:0] ki6=212;
reg signed [w1-1:0] ka7=-129;	reg signed [w1-1:0] kb7=-237;	reg signed [w1-1:0] kc7=254;	reg signed [w1-1:0] kd7=-111;	reg signed [w1-1:0] ke7=-74;	reg signed [w1-1:0] kf7=-208;	reg signed [w1-1:0] kg7=285;	reg signed [w1-1:0] kh7=-118;	reg signed [w1-1:0] ki7=-167;
reg signed [w1-1:0] ka8=109;	reg signed [w1-1:0] kb8=90;	reg signed [w1-1:0] kc8=-363;	reg signed [w1-1:0] kd8=-182;	reg signed [w1-1:0] ke8=-218;	reg signed [w1-1:0] kf8=-41;	reg signed [w1-1:0] kg8=25;	reg signed [w1-1:0] kh8=-41;	reg signed [w1-1:0] ki8=414;


reg signed [w4-1:0] delta1=36;	reg signed [w4-1:0] mu1=-321;	reg signed [w4-1:0] beta1=-5558;
reg signed [w4-1:0] delta2=41;	reg signed [w4-1:0] mu2=323;	reg signed [w4-1:0] beta2=-11873;
reg signed [w4-1:0] delta3=47;	reg signed [w4-1:0] mu3=137;	reg signed [w4-1:0] beta3=56083;
reg signed [w4-1:0] delta4=44;	reg signed [w4-1:0] mu4=-24;	reg signed [w4-1:0] beta4=86292;
reg signed [w4-1:0] delta5=48;	reg signed [w4-1:0] mu5=86;	reg signed [w4-1:0] beta5=-33672;
reg signed [w4-1:0] delta6=18;	reg signed [w4-1:0] mu6=996;	reg signed [w4-1:0] beta6=60113;
reg signed [w4-1:0] delta7=36;	reg signed [w4-1:0] mu7=-48;	reg signed [w4-1:0] beta7=-63190;
reg signed [w4-1:0] delta8=40;	reg signed [w4-1:0] mu8=182;	reg signed [w4-1:0] beta8=-53799;


reg signed [w5-1:0] ka9=101;	reg signed [w5-1:0] kb9=110;	reg signed [w5-1:0] kc9=152;	reg signed [w5-1:0] kd9=-43;	reg signed [w5-1:0] ke9=-94;	reg signed [w5-1:0] kf9=93;	reg signed [w5-1:0] kg9=62;	reg signed [w5-1:0] kh9=75;	reg signed [w5-1:0] ki9=-39;
reg signed [w5-1:0] ka10=-65;	reg signed [w5-1:0] kb10=-20;	reg signed [w5-1:0] kc10=107;	reg signed [w5-1:0] kd10=-14;	reg signed [w5-1:0] ke10=-124;	reg signed [w5-1:0] kf10=-57;	reg signed [w5-1:0] kg10=-105;	reg signed [w5-1:0] kh10=12;	reg signed [w5-1:0] ki10=-68;
reg signed [w5-1:0] ka11=-165;	reg signed [w5-1:0] kb11=-95;	reg signed [w5-1:0] kc11=-145;	reg signed [w5-1:0] kd11=66;	reg signed [w5-1:0] ke11=30;	reg signed [w5-1:0] kf11=5;	reg signed [w5-1:0] kg11=-87;	reg signed [w5-1:0] kh11=147;	reg signed [w5-1:0] ki11=197;
reg signed [w5-1:0] ka12=36;	reg signed [w5-1:0] kb12=-78;	reg signed [w5-1:0] kc12=-116;	reg signed [w5-1:0] kd12=-175;	reg signed [w5-1:0] ke12=-28;	reg signed [w5-1:0] kf12=5;	reg signed [w5-1:0] kg12=-138;	reg signed [w5-1:0] kh12=106;	reg signed [w5-1:0] ki12=165;
reg signed [w5-1:0] ka13=114;	reg signed [w5-1:0] kb13=-140;	reg signed [w5-1:0] kc13=-147;	reg signed [w5-1:0] kd13=-39;	reg signed [w5-1:0] ke13=-119;	reg signed [w5-1:0] kf13=-11;	reg signed [w5-1:0] kg13=117;	reg signed [w5-1:0] kh13=156;	reg signed [w5-1:0] ki13=-48;
reg signed [w5-1:0] ka14=-187;	reg signed [w5-1:0] kb14=-107;	reg signed [w5-1:0] kc14=148;	reg signed [w5-1:0] kd14=-147;	reg signed [w5-1:0] ke14=64;	reg signed [w5-1:0] kf14=67;	reg signed [w5-1:0] kg14=20;	reg signed [w5-1:0] kh14=-27;	reg signed [w5-1:0] ki14=-50;
reg signed [w5-1:0] ka15=26;	reg signed [w5-1:0] kb15=128;	reg signed [w5-1:0] kc15=-112;	reg signed [w5-1:0] kd15=86;	reg signed [w5-1:0] ke15=-37;	reg signed [w5-1:0] kf15=65;	reg signed [w5-1:0] kg15=-5;	reg signed [w5-1:0] kh15=-40;	reg signed [w5-1:0] ki15=-79;
reg signed [w5-1:0] ka16=-5;	reg signed [w5-1:0] kb16=56;	reg signed [w5-1:0] kc16=78;	reg signed [w5-1:0] kd16=-50;	reg signed [w5-1:0] ke16=180;	reg signed [w5-1:0] kf16=128;	reg signed [w5-1:0] kg16=1;	reg signed [w5-1:0] kh16=132;	reg signed [w5-1:0] ki16=-153;
reg signed [w5-1:0] ka17=41;	reg signed [w5-1:0] kb17=-39;	reg signed [w5-1:0] kc17=176;	reg signed [w5-1:0] kd17=153;	reg signed [w5-1:0] ke17=-121;	reg signed [w5-1:0] kf17=66;	reg signed [w5-1:0] kg17=0;	reg signed [w5-1:0] kh17=50;	reg signed [w5-1:0] ki17=-43;
reg signed [w5-1:0] ka18=26;	reg signed [w5-1:0] kb18=16;	reg signed [w5-1:0] kc18=12;	reg signed [w5-1:0] kd18=44;	reg signed [w5-1:0] ke18=-36;	reg signed [w5-1:0] kf18=66;	reg signed [w5-1:0] kg18=145;	reg signed [w5-1:0] kh18=127;	reg signed [w5-1:0] ki18=47;
reg signed [w5-1:0] ka19=155;	reg signed [w5-1:0] kb19=11;	reg signed [w5-1:0] kc19=90;	reg signed [w5-1:0] kd19=-6;	reg signed [w5-1:0] ke19=2;	reg signed [w5-1:0] kf19=-25;	reg signed [w5-1:0] kg19=87;	reg signed [w5-1:0] kh19=3;	reg signed [w5-1:0] ki19=201;
reg signed [w5-1:0] ka20=167;	reg signed [w5-1:0] kb20=166;	reg signed [w5-1:0] kc20=70;	reg signed [w5-1:0] kd20=-104;	reg signed [w5-1:0] ke20=78;	reg signed [w5-1:0] kf20=116;	reg signed [w5-1:0] kg20=-61;	reg signed [w5-1:0] kh20=98;	reg signed [w5-1:0] ki20=24;
reg signed [w5-1:0] ka21=153;	reg signed [w5-1:0] kb21=51;	reg signed [w5-1:0] kc21=-10;	reg signed [w5-1:0] kd21=-104;	reg signed [w5-1:0] ke21=-46;	reg signed [w5-1:0] kf21=124;	reg signed [w5-1:0] kg21=30;	reg signed [w5-1:0] kh21=14;	reg signed [w5-1:0] ki21=49;
reg signed [w5-1:0] ka22=144;	reg signed [w5-1:0] kb22=-200;	reg signed [w5-1:0] kc22=138;	reg signed [w5-1:0] kd22=129;	reg signed [w5-1:0] ke22=-40;	reg signed [w5-1:0] kf22=27;	reg signed [w5-1:0] kg22=39;	reg signed [w5-1:0] kh22=-128;	reg signed [w5-1:0] ki22=171;
reg signed [w5-1:0] ka23=25;	reg signed [w5-1:0] kb23=144;	reg signed [w5-1:0] kc23=-39;	reg signed [w5-1:0] kd23=-23;	reg signed [w5-1:0] ke23=7;	reg signed [w5-1:0] kf23=114;	reg signed [w5-1:0] kg23=-130;	reg signed [w5-1:0] kh23=-111;	reg signed [w5-1:0] ki23=-1;
reg signed [w5-1:0] ka24=-30;	reg signed [w5-1:0] kb24=-93;	reg signed [w5-1:0] kc24=11;	reg signed [w5-1:0] kd24=-38;	reg signed [w5-1:0] ke24=-39;	reg signed [w5-1:0] kf24=-25;	reg signed [w5-1:0] kg24=-114;	reg signed [w5-1:0] kh24=-9;	reg signed [w5-1:0] ki24=106;
reg signed [w5-1:0] ka25=-34;	reg signed [w5-1:0] kb25=-44;	reg signed [w5-1:0] kc25=-6;	reg signed [w5-1:0] kd25=77;	reg signed [w5-1:0] ke25=-32;	reg signed [w5-1:0] kf25=6;	reg signed [w5-1:0] kg25=-68;	reg signed [w5-1:0] kh25=124;	reg signed [w5-1:0] ki25=-97;
reg signed [w5-1:0] ka26=-152;	reg signed [w5-1:0] kb26=-154;	reg signed [w5-1:0] kc26=28;	reg signed [w5-1:0] kd26=5;	reg signed [w5-1:0] ke26=-144;	reg signed [w5-1:0] kf26=12;	reg signed [w5-1:0] kg26=166;	reg signed [w5-1:0] kh26=-153;	reg signed [w5-1:0] ki26=-36;
reg signed [w5-1:0] ka27=155;	reg signed [w5-1:0] kb27=148;	reg signed [w5-1:0] kc27=-17;	reg signed [w5-1:0] kd27=12;	reg signed [w5-1:0] ke27=-107;	reg signed [w5-1:0] kf27=83;	reg signed [w5-1:0] kg27=-7;	reg signed [w5-1:0] kh27=69;	reg signed [w5-1:0] ki27=74;
reg signed [w5-1:0] ka28=-87;	reg signed [w5-1:0] kb28=-58;	reg signed [w5-1:0] kc28=96;	reg signed [w5-1:0] kd28=51;	reg signed [w5-1:0] ke28=18;	reg signed [w5-1:0] kf28=105;	reg signed [w5-1:0] kg28=-81;	reg signed [w5-1:0] kh28=142;	reg signed [w5-1:0] ki28=-14;
reg signed [w5-1:0] ka29=46;	reg signed [w5-1:0] kb29=54;	reg signed [w5-1:0] kc29=11;	reg signed [w5-1:0] kd29=148;	reg signed [w5-1:0] ke29=-150;	reg signed [w5-1:0] kf29=-143;	reg signed [w5-1:0] kg29=-127;	reg signed [w5-1:0] kh29=-6;	reg signed [w5-1:0] ki29=69;
reg signed [w5-1:0] ka30=58;	reg signed [w5-1:0] kb30=-33;	reg signed [w5-1:0] kc30=-104;	reg signed [w5-1:0] kd30=192;	reg signed [w5-1:0] ke30=62;	reg signed [w5-1:0] kf30=78;	reg signed [w5-1:0] kg30=97;	reg signed [w5-1:0] kh30=63;	reg signed [w5-1:0] ki30=219;
reg signed [w5-1:0] ka31=-27;	reg signed [w5-1:0] kb31=-104;	reg signed [w5-1:0] kc31=38;	reg signed [w5-1:0] kd31=28;	reg signed [w5-1:0] ke31=30;	reg signed [w5-1:0] kf31=-136;	reg signed [w5-1:0] kg31=36;	reg signed [w5-1:0] kh31=-117;	reg signed [w5-1:0] ki31=-104;
reg signed [w5-1:0] ka32=115;	reg signed [w5-1:0] kb32=52;	reg signed [w5-1:0] kc32=183;	reg signed [w5-1:0] kd32=-65;	reg signed [w5-1:0] ke32=-65;	reg signed [w5-1:0] kf32=52;	reg signed [w5-1:0] kg32=-89;	reg signed [w5-1:0] kh32=-63;	reg signed [w5-1:0] ki32=-154;
reg signed [w5-1:0] ka33=-116;	reg signed [w5-1:0] kb33=12;	reg signed [w5-1:0] kc33=125;	reg signed [w5-1:0] kd33=-36;	reg signed [w5-1:0] ke33=-87;	reg signed [w5-1:0] kf33=107;	reg signed [w5-1:0] kg33=177;	reg signed [w5-1:0] kh33=-8;	reg signed [w5-1:0] ki33=12;
reg signed [w5-1:0] ka34=-115;	reg signed [w5-1:0] kb34=69;	reg signed [w5-1:0] kc34=-132;	reg signed [w5-1:0] kd34=4;	reg signed [w5-1:0] ke34=-124;	reg signed [w5-1:0] kf34=-84;	reg signed [w5-1:0] kg34=-103;	reg signed [w5-1:0] kh34=-142;	reg signed [w5-1:0] ki34=-7;
reg signed [w5-1:0] ka35=137;	reg signed [w5-1:0] kb35=-46;	reg signed [w5-1:0] kc35=-192;	reg signed [w5-1:0] kd35=128;	reg signed [w5-1:0] ke35=0;	reg signed [w5-1:0] kf35=5;	reg signed [w5-1:0] kg35=-34;	reg signed [w5-1:0] kh35=102;	reg signed [w5-1:0] ki35=52;
reg signed [w5-1:0] ka36=-20;	reg signed [w5-1:0] kb36=-97;	reg signed [w5-1:0] kc36=-133;	reg signed [w5-1:0] kd36=31;	reg signed [w5-1:0] ke36=46;	reg signed [w5-1:0] kf36=172;	reg signed [w5-1:0] kg36=-32;	reg signed [w5-1:0] kh36=-130;	reg signed [w5-1:0] ki36=-2;
reg signed [w5-1:0] ka37=-136;	reg signed [w5-1:0] kb37=-144;	reg signed [w5-1:0] kc37=139;	reg signed [w5-1:0] kd37=155;	reg signed [w5-1:0] ke37=-105;	reg signed [w5-1:0] kf37=-145;	reg signed [w5-1:0] kg37=-151;	reg signed [w5-1:0] kh37=81;	reg signed [w5-1:0] ki37=42;
reg signed [w5-1:0] ka38=129;	reg signed [w5-1:0] kb38=-44;	reg signed [w5-1:0] kc38=-158;	reg signed [w5-1:0] kd38=197;	reg signed [w5-1:0] ke38=140;	reg signed [w5-1:0] kf38=-67;	reg signed [w5-1:0] kg38=202;	reg signed [w5-1:0] kh38=-3;	reg signed [w5-1:0] ki38=55;
reg signed [w5-1:0] ka39=159;	reg signed [w5-1:0] kb39=181;	reg signed [w5-1:0] kc39=-46;	reg signed [w5-1:0] kd39=148;	reg signed [w5-1:0] ke39=-10;	reg signed [w5-1:0] kf39=-99;	reg signed [w5-1:0] kg39=24;	reg signed [w5-1:0] kh39=-128;	reg signed [w5-1:0] ki39=152;
reg signed [w5-1:0] ka40=-103;	reg signed [w5-1:0] kb40=-120;	reg signed [w5-1:0] kc40=138;	reg signed [w5-1:0] kd40=-145;	reg signed [w5-1:0] ke40=-97;	reg signed [w5-1:0] kf40=-60;	reg signed [w5-1:0] kg40=-100;	reg signed [w5-1:0] kh40=111;	reg signed [w5-1:0] ki40=-66;
reg signed [w5-1:0] ka41=24;	reg signed [w5-1:0] kb41=113;	reg signed [w5-1:0] kc41=-59;	reg signed [w5-1:0] kd41=6;	reg signed [w5-1:0] ke41=-80;	reg signed [w5-1:0] kf41=33;	reg signed [w5-1:0] kg41=-99;	reg signed [w5-1:0] kh41=107;	reg signed [w5-1:0] ki41=-89;
reg signed [w5-1:0] ka42=-191;	reg signed [w5-1:0] kb42=38;	reg signed [w5-1:0] kc42=226;	reg signed [w5-1:0] kd42=153;	reg signed [w5-1:0] ke42=78;	reg signed [w5-1:0] kf42=55;	reg signed [w5-1:0] kg42=-1;	reg signed [w5-1:0] kh42=132;	reg signed [w5-1:0] ki42=177;
reg signed [w5-1:0] ka43=173;	reg signed [w5-1:0] kb43=-81;	reg signed [w5-1:0] kc43=174;	reg signed [w5-1:0] kd43=99;	reg signed [w5-1:0] ke43=-171;	reg signed [w5-1:0] kf43=81;	reg signed [w5-1:0] kg43=-68;	reg signed [w5-1:0] kh43=47;	reg signed [w5-1:0] ki43=26;
reg signed [w5-1:0] ka44=-109;	reg signed [w5-1:0] kb44=-19;	reg signed [w5-1:0] kc44=-106;	reg signed [w5-1:0] kd44=-26;	reg signed [w5-1:0] ke44=94;	reg signed [w5-1:0] kf44=6;	reg signed [w5-1:0] kg44=27;	reg signed [w5-1:0] kh44=86;	reg signed [w5-1:0] ki44=32;
reg signed [w5-1:0] ka45=0;	reg signed [w5-1:0] kb45=-109;	reg signed [w5-1:0] kc45=4;	reg signed [w5-1:0] kd45=-123;	reg signed [w5-1:0] ke45=-73;	reg signed [w5-1:0] kf45=155;	reg signed [w5-1:0] kg45=-161;	reg signed [w5-1:0] kh45=13;	reg signed [w5-1:0] ki45=92;
reg signed [w5-1:0] ka46=131;	reg signed [w5-1:0] kb46=144;	reg signed [w5-1:0] kc46=126;	reg signed [w5-1:0] kd46=-173;	reg signed [w5-1:0] ke46=-131;	reg signed [w5-1:0] kf46=-149;	reg signed [w5-1:0] kg46=66;	reg signed [w5-1:0] kh46=144;	reg signed [w5-1:0] ki46=53;
reg signed [w5-1:0] ka47=-118;	reg signed [w5-1:0] kb47=-84;	reg signed [w5-1:0] kc47=-70;	reg signed [w5-1:0] kd47=-161;	reg signed [w5-1:0] ke47=-39;	reg signed [w5-1:0] kf47=54;	reg signed [w5-1:0] kg47=-88;	reg signed [w5-1:0] kh47=-69;	reg signed [w5-1:0] ki47=158;
reg signed [w5-1:0] ka48=-160;	reg signed [w5-1:0] kb48=65;	reg signed [w5-1:0] kc48=-105;	reg signed [w5-1:0] kd48=-41;	reg signed [w5-1:0] ke48=80;	reg signed [w5-1:0] kf48=21;	reg signed [w5-1:0] kg48=34;	reg signed [w5-1:0] kh48=46;	reg signed [w5-1:0] ki48=113;
reg signed [w5-1:0] ka49=-241;	reg signed [w5-1:0] kb49=-84;	reg signed [w5-1:0] kc49=-215;	reg signed [w5-1:0] kd49=-94;	reg signed [w5-1:0] ke49=-109;	reg signed [w5-1:0] kf49=-184;	reg signed [w5-1:0] kg49=-69;	reg signed [w5-1:0] kh49=180;	reg signed [w5-1:0] ki49=123;
reg signed [w5-1:0] ka50=-6;	reg signed [w5-1:0] kb50=26;	reg signed [w5-1:0] kc50=185;	reg signed [w5-1:0] kd50=-65;	reg signed [w5-1:0] ke50=125;	reg signed [w5-1:0] kf50=-67;	reg signed [w5-1:0] kg50=-77;	reg signed [w5-1:0] kh50=89;	reg signed [w5-1:0] ki50=-18;
reg signed [w5-1:0] ka51=-126;	reg signed [w5-1:0] kb51=92;	reg signed [w5-1:0] kc51=78;	reg signed [w5-1:0] kd51=102;	reg signed [w5-1:0] ke51=-135;	reg signed [w5-1:0] kf51=-86;	reg signed [w5-1:0] kg51=185;	reg signed [w5-1:0] kh51=-122;	reg signed [w5-1:0] ki51=34;
reg signed [w5-1:0] ka52=-29;	reg signed [w5-1:0] kb52=82;	reg signed [w5-1:0] kc52=-45;	reg signed [w5-1:0] kd52=29;	reg signed [w5-1:0] ke52=-27;	reg signed [w5-1:0] kf52=-17;	reg signed [w5-1:0] kg52=-142;	reg signed [w5-1:0] kh52=-21;	reg signed [w5-1:0] ki52=50;
reg signed [w5-1:0] ka53=50;	reg signed [w5-1:0] kb53=-117;	reg signed [w5-1:0] kc53=57;	reg signed [w5-1:0] kd53=79;	reg signed [w5-1:0] ke53=-2;	reg signed [w5-1:0] kf53=-3;	reg signed [w5-1:0] kg53=-96;	reg signed [w5-1:0] kh53=161;	reg signed [w5-1:0] ki53=-47;
reg signed [w5-1:0] ka54=154;	reg signed [w5-1:0] kb54=40;	reg signed [w5-1:0] kc54=61;	reg signed [w5-1:0] kd54=-81;	reg signed [w5-1:0] ke54=43;	reg signed [w5-1:0] kf54=179;	reg signed [w5-1:0] kg54=-192;	reg signed [w5-1:0] kh54=54;	reg signed [w5-1:0] ki54=-92;
reg signed [w5-1:0] ka55=173;	reg signed [w5-1:0] kb55=152;	reg signed [w5-1:0] kc55=53;	reg signed [w5-1:0] kd55=154;	reg signed [w5-1:0] ke55=187;	reg signed [w5-1:0] kf55=98;	reg signed [w5-1:0] kg55=21;	reg signed [w5-1:0] kh55=144;	reg signed [w5-1:0] ki55=148;
reg signed [w5-1:0] ka56=88;	reg signed [w5-1:0] kb56=112;	reg signed [w5-1:0] kc56=-154;	reg signed [w5-1:0] kd56=150;	reg signed [w5-1:0] ke56=141;	reg signed [w5-1:0] kf56=114;	reg signed [w5-1:0] kg56=-52;	reg signed [w5-1:0] kh56=-28;	reg signed [w5-1:0] ki56=66;
reg signed [w5-1:0] ka57=214;	reg signed [w5-1:0] kb57=90;	reg signed [w5-1:0] kc57=-62;	reg signed [w5-1:0] kd57=14;	reg signed [w5-1:0] ke57=144;	reg signed [w5-1:0] kf57=-22;	reg signed [w5-1:0] kg57=-128;	reg signed [w5-1:0] kh57=-58;	reg signed [w5-1:0] ki57=-62;
reg signed [w5-1:0] ka58=-145;	reg signed [w5-1:0] kb58=14;	reg signed [w5-1:0] kc58=89;	reg signed [w5-1:0] kd58=65;	reg signed [w5-1:0] ke58=-16;	reg signed [w5-1:0] kf58=119;	reg signed [w5-1:0] kg58=197;	reg signed [w5-1:0] kh58=241;	reg signed [w5-1:0] ki58=107;
reg signed [w5-1:0] ka59=87;	reg signed [w5-1:0] kb59=180;	reg signed [w5-1:0] kc59=-2;	reg signed [w5-1:0] kd59=10;	reg signed [w5-1:0] ke59=-22;	reg signed [w5-1:0] kf59=57;	reg signed [w5-1:0] kg59=111;	reg signed [w5-1:0] kh59=8;	reg signed [w5-1:0] ki59=-87;
reg signed [w5-1:0] ka60=-58;	reg signed [w5-1:0] kb60=164;	reg signed [w5-1:0] kc60=-86;	reg signed [w5-1:0] kd60=-47;	reg signed [w5-1:0] ke60=58;	reg signed [w5-1:0] kf60=41;	reg signed [w5-1:0] kg60=56;	reg signed [w5-1:0] kh60=20;	reg signed [w5-1:0] ki60=187;
reg signed [w5-1:0] ka61=186;	reg signed [w5-1:0] kb61=-103;	reg signed [w5-1:0] kc61=-150;	reg signed [w5-1:0] kd61=-7;	reg signed [w5-1:0] ke61=95;	reg signed [w5-1:0] kf61=-36;	reg signed [w5-1:0] kg61=-37;	reg signed [w5-1:0] kh61=39;	reg signed [w5-1:0] ki61=-9;
reg signed [w5-1:0] ka62=68;	reg signed [w5-1:0] kb62=-146;	reg signed [w5-1:0] kc62=7;	reg signed [w5-1:0] kd62=132;	reg signed [w5-1:0] ke62=10;	reg signed [w5-1:0] kf62=-83;	reg signed [w5-1:0] kg62=52;	reg signed [w5-1:0] kh62=30;	reg signed [w5-1:0] ki62=-56;
reg signed [w5-1:0] ka63=150;	reg signed [w5-1:0] kb63=11;	reg signed [w5-1:0] kc63=43;	reg signed [w5-1:0] kd63=3;	reg signed [w5-1:0] ke63=77;	reg signed [w5-1:0] kf63=21;	reg signed [w5-1:0] kg63=158;	reg signed [w5-1:0] kh63=163;	reg signed [w5-1:0] ki63=31;
reg signed [w5-1:0] ka64=-66;	reg signed [w5-1:0] kb64=50;	reg signed [w5-1:0] kc64=-103;	reg signed [w5-1:0] kd64=129;	reg signed [w5-1:0] ke64=9;	reg signed [w5-1:0] kf64=59;	reg signed [w5-1:0] kg64=127;	reg signed [w5-1:0] kh64=16;	reg signed [w5-1:0] ki64=73;
reg signed [w5-1:0] ka65=8;	reg signed [w5-1:0] kb65=-91;	reg signed [w5-1:0] kc65=72;	reg signed [w5-1:0] kd65=-173;	reg signed [w5-1:0] ke65=-28;	reg signed [w5-1:0] kf65=105;	reg signed [w5-1:0] kg65=-132;	reg signed [w5-1:0] kh65=137;	reg signed [w5-1:0] ki65=-99;
reg signed [w5-1:0] ka66=-146;	reg signed [w5-1:0] kb66=55;	reg signed [w5-1:0] kc66=-72;	reg signed [w5-1:0] kd66=-102;	reg signed [w5-1:0] ke66=-83;	reg signed [w5-1:0] kf66=-86;	reg signed [w5-1:0] kg66=-7;	reg signed [w5-1:0] kh66=-78;	reg signed [w5-1:0] ki66=-107;
reg signed [w5-1:0] ka67=35;	reg signed [w5-1:0] kb67=139;	reg signed [w5-1:0] kc67=80;	reg signed [w5-1:0] kd67=-32;	reg signed [w5-1:0] ke67=122;	reg signed [w5-1:0] kf67=-49;	reg signed [w5-1:0] kg67=153;	reg signed [w5-1:0] kh67=152;	reg signed [w5-1:0] ki67=186;
reg signed [w5-1:0] ka68=194;	reg signed [w5-1:0] kb68=-61;	reg signed [w5-1:0] kc68=-59;	reg signed [w5-1:0] kd68=181;	reg signed [w5-1:0] ke68=-19;	reg signed [w5-1:0] kf68=-8;	reg signed [w5-1:0] kg68=-84;	reg signed [w5-1:0] kh68=82;	reg signed [w5-1:0] ki68=151;
reg signed [w5-1:0] ka69=-27;	reg signed [w5-1:0] kb69=-63;	reg signed [w5-1:0] kc69=57;	reg signed [w5-1:0] kd69=-148;	reg signed [w5-1:0] ke69=-77;	reg signed [w5-1:0] kf69=4;	reg signed [w5-1:0] kg69=191;	reg signed [w5-1:0] kh69=-24;	reg signed [w5-1:0] ki69=-49;
reg signed [w5-1:0] ka70=73;	reg signed [w5-1:0] kb70=113;	reg signed [w5-1:0] kc70=-34;	reg signed [w5-1:0] kd70=-122;	reg signed [w5-1:0] ke70=32;	reg signed [w5-1:0] kf70=97;	reg signed [w5-1:0] kg70=28;	reg signed [w5-1:0] kh70=128;	reg signed [w5-1:0] ki70=-78;
reg signed [w5-1:0] ka71=-10;	reg signed [w5-1:0] kb71=-129;	reg signed [w5-1:0] kc71=89;	reg signed [w5-1:0] kd71=-9;	reg signed [w5-1:0] ke71=-92;	reg signed [w5-1:0] kf71=-137;	reg signed [w5-1:0] kg71=-181;	reg signed [w5-1:0] kh71=-86;	reg signed [w5-1:0] ki71=128;
reg signed [w5-1:0] ka72=-191;	reg signed [w5-1:0] kb72=145;	reg signed [w5-1:0] kc72=6;	reg signed [w5-1:0] kd72=-68;	reg signed [w5-1:0] ke72=-57;	reg signed [w5-1:0] kf72=-10;	reg signed [w5-1:0] kg72=34;	reg signed [w5-1:0] kh72=165;	reg signed [w5-1:0] ki72=129;
reg signed [w5-1:0] ka73=17;	reg signed [w5-1:0] kb73=-72;	reg signed [w5-1:0] kc73=75;	reg signed [w5-1:0] kd73=-77;	reg signed [w5-1:0] ke73=68;	reg signed [w5-1:0] kf73=48;	reg signed [w5-1:0] kg73=74;	reg signed [w5-1:0] kh73=-1;	reg signed [w5-1:0] ki73=-74;
reg signed [w5-1:0] ka74=89;	reg signed [w5-1:0] kb74=132;	reg signed [w5-1:0] kc74=38;	reg signed [w5-1:0] kd74=115;	reg signed [w5-1:0] ke74=-17;	reg signed [w5-1:0] kf74=186;	reg signed [w5-1:0] kg74=-96;	reg signed [w5-1:0] kh74=59;	reg signed [w5-1:0] ki74=-49;
reg signed [w5-1:0] ka75=74;	reg signed [w5-1:0] kb75=-48;	reg signed [w5-1:0] kc75=2;	reg signed [w5-1:0] kd75=-66;	reg signed [w5-1:0] ke75=79;	reg signed [w5-1:0] kf75=69;	reg signed [w5-1:0] kg75=-30;	reg signed [w5-1:0] kh75=127;	reg signed [w5-1:0] ki75=131;
reg signed [w5-1:0] ka76=121;	reg signed [w5-1:0] kb76=-52;	reg signed [w5-1:0] kc76=-100;	reg signed [w5-1:0] kd76=104;	reg signed [w5-1:0] ke76=-99;	reg signed [w5-1:0] kf76=104;	reg signed [w5-1:0] kg76=2;	reg signed [w5-1:0] kh76=76;	reg signed [w5-1:0] ki76=145;
reg signed [w5-1:0] ka77=34;	reg signed [w5-1:0] kb77=198;	reg signed [w5-1:0] kc77=169;	reg signed [w5-1:0] kd77=-64;	reg signed [w5-1:0] ke77=84;	reg signed [w5-1:0] kf77=147;	reg signed [w5-1:0] kg77=-148;	reg signed [w5-1:0] kh77=65;	reg signed [w5-1:0] ki77=101;
reg signed [w5-1:0] ka78=21;	reg signed [w5-1:0] kb78=-36;	reg signed [w5-1:0] kc78=-186;	reg signed [w5-1:0] kd78=121;	reg signed [w5-1:0] ke78=-56;	reg signed [w5-1:0] kf78=127;	reg signed [w5-1:0] kg78=-182;	reg signed [w5-1:0] kh78=-201;	reg signed [w5-1:0] ki78=-202;
reg signed [w5-1:0] ka79=106;	reg signed [w5-1:0] kb79=-183;	reg signed [w5-1:0] kc79=124;	reg signed [w5-1:0] kd79=28;	reg signed [w5-1:0] ke79=96;	reg signed [w5-1:0] kf79=-78;	reg signed [w5-1:0] kg79=-137;	reg signed [w5-1:0] kh79=-46;	reg signed [w5-1:0] ki79=89;
reg signed [w5-1:0] ka80=-61;	reg signed [w5-1:0] kb80=53;	reg signed [w5-1:0] kc80=63;	reg signed [w5-1:0] kd80=196;	reg signed [w5-1:0] ke80=158;	reg signed [w5-1:0] kf80=69;	reg signed [w5-1:0] kg80=158;	reg signed [w5-1:0] kh80=107;	reg signed [w5-1:0] ki80=-127;
reg signed [w5-1:0] ka81=137;	reg signed [w5-1:0] kb81=-57;	reg signed [w5-1:0] kc81=-55;	reg signed [w5-1:0] kd81=20;	reg signed [w5-1:0] ke81=-131;	reg signed [w5-1:0] kf81=-127;	reg signed [w5-1:0] kg81=226;	reg signed [w5-1:0] kh81=63;	reg signed [w5-1:0] ki81=124;
reg signed [w5-1:0] ka82=-3;	reg signed [w5-1:0] kb82=60;	reg signed [w5-1:0] kc82=101;	reg signed [w5-1:0] kd82=104;	reg signed [w5-1:0] ke82=94;	reg signed [w5-1:0] kf82=-25;	reg signed [w5-1:0] kg82=-35;	reg signed [w5-1:0] kh82=-46;	reg signed [w5-1:0] ki82=-103;
reg signed [w5-1:0] ka83=-2;	reg signed [w5-1:0] kb83=54;	reg signed [w5-1:0] kc83=61;	reg signed [w5-1:0] kd83=-111;	reg signed [w5-1:0] ke83=4;	reg signed [w5-1:0] kf83=90;	reg signed [w5-1:0] kg83=-98;	reg signed [w5-1:0] kh83=-9;	reg signed [w5-1:0] ki83=-194;
reg signed [w5-1:0] ka84=80;	reg signed [w5-1:0] kb84=142;	reg signed [w5-1:0] kc84=-25;	reg signed [w5-1:0] kd84=-19;	reg signed [w5-1:0] ke84=-123;	reg signed [w5-1:0] kf84=81;	reg signed [w5-1:0] kg84=-11;	reg signed [w5-1:0] kh84=-197;	reg signed [w5-1:0] ki84=-24;
reg signed [w5-1:0] ka85=-27;	reg signed [w5-1:0] kb85=31;	reg signed [w5-1:0] kc85=5;	reg signed [w5-1:0] kd85=-131;	reg signed [w5-1:0] ke85=37;	reg signed [w5-1:0] kf85=177;	reg signed [w5-1:0] kg85=-104;	reg signed [w5-1:0] kh85=-14;	reg signed [w5-1:0] ki85=-18;
reg signed [w5-1:0] ka86=-17;	reg signed [w5-1:0] kb86=-3;	reg signed [w5-1:0] kc86=124;	reg signed [w5-1:0] kd86=-109;	reg signed [w5-1:0] ke86=-119;	reg signed [w5-1:0] kf86=142;	reg signed [w5-1:0] kg86=49;	reg signed [w5-1:0] kh86=-34;	reg signed [w5-1:0] ki86=24;
reg signed [w5-1:0] ka87=70;	reg signed [w5-1:0] kb87=-75;	reg signed [w5-1:0] kc87=34;	reg signed [w5-1:0] kd87=67;	reg signed [w5-1:0] ke87=148;	reg signed [w5-1:0] kf87=150;	reg signed [w5-1:0] kg87=-46;	reg signed [w5-1:0] kh87=234;	reg signed [w5-1:0] ki87=-29;
reg signed [w5-1:0] ka88=1;	reg signed [w5-1:0] kb88=81;	reg signed [w5-1:0] kc88=134;	reg signed [w5-1:0] kd88=-141;	reg signed [w5-1:0] ke88=-77;	reg signed [w5-1:0] kf88=58;	reg signed [w5-1:0] kg88=-224;	reg signed [w5-1:0] kh88=-203;	reg signed [w5-1:0] ki88=8;
reg signed [w5-1:0] ka89=-81;	reg signed [w5-1:0] kb89=5;	reg signed [w5-1:0] kc89=-63;	reg signed [w5-1:0] kd89=38;	reg signed [w5-1:0] ke89=-39;	reg signed [w5-1:0] kf89=105;	reg signed [w5-1:0] kg89=-34;	reg signed [w5-1:0] kh89=-41;	reg signed [w5-1:0] ki89=-71;
reg signed [w5-1:0] ka90=160;	reg signed [w5-1:0] kb90=-83;	reg signed [w5-1:0] kc90=-79;	reg signed [w5-1:0] kd90=166;	reg signed [w5-1:0] ke90=-86;	reg signed [w5-1:0] kf90=-50;	reg signed [w5-1:0] kg90=-79;	reg signed [w5-1:0] kh90=-79;	reg signed [w5-1:0] ki90=148;
reg signed [w5-1:0] ka91=43;	reg signed [w5-1:0] kb91=157;	reg signed [w5-1:0] kc91=-78;	reg signed [w5-1:0] kd91=-137;	reg signed [w5-1:0] ke91=-135;	reg signed [w5-1:0] kf91=-17;	reg signed [w5-1:0] kg91=64;	reg signed [w5-1:0] kh91=106;	reg signed [w5-1:0] ki91=-69;
reg signed [w5-1:0] ka92=6;	reg signed [w5-1:0] kb92=56;	reg signed [w5-1:0] kc92=-12;	reg signed [w5-1:0] kd92=-85;	reg signed [w5-1:0] ke92=-137;	reg signed [w5-1:0] kf92=-83;	reg signed [w5-1:0] kg92=-142;	reg signed [w5-1:0] kh92=-88;	reg signed [w5-1:0] ki92=-80;
reg signed [w5-1:0] ka93=87;	reg signed [w5-1:0] kb93=159;	reg signed [w5-1:0] kc93=-155;	reg signed [w5-1:0] kd93=-161;	reg signed [w5-1:0] ke93=-147;	reg signed [w5-1:0] kf93=39;	reg signed [w5-1:0] kg93=99;	reg signed [w5-1:0] kh93=-108;	reg signed [w5-1:0] ki93=64;
reg signed [w5-1:0] ka94=107;	reg signed [w5-1:0] kb94=8;	reg signed [w5-1:0] kc94=-45;	reg signed [w5-1:0] kd94=-109;	reg signed [w5-1:0] ke94=-136;	reg signed [w5-1:0] kf94=126;	reg signed [w5-1:0] kg94=146;	reg signed [w5-1:0] kh94=-81;	reg signed [w5-1:0] ki94=-155;
reg signed [w5-1:0] ka95=-60;	reg signed [w5-1:0] kb95=-149;	reg signed [w5-1:0] kc95=-56;	reg signed [w5-1:0] kd95=66;	reg signed [w5-1:0] ke95=113;	reg signed [w5-1:0] kf95=-65;	reg signed [w5-1:0] kg95=126;	reg signed [w5-1:0] kh95=-139;	reg signed [w5-1:0] ki95=162;
reg signed [w5-1:0] ka96=56;	reg signed [w5-1:0] kb96=-105;	reg signed [w5-1:0] kc96=-176;	reg signed [w5-1:0] kd96=4;	reg signed [w5-1:0] ke96=102;	reg signed [w5-1:0] kf96=-158;	reg signed [w5-1:0] kg96=83;	reg signed [w5-1:0] kh96=5;	reg signed [w5-1:0] ki96=-69;
reg signed [w5-1:0] ka97=-171;	reg signed [w5-1:0] kb97=38;	reg signed [w5-1:0] kc97=76;	reg signed [w5-1:0] kd97=41;	reg signed [w5-1:0] ke97=7;	reg signed [w5-1:0] kf97=-60;	reg signed [w5-1:0] kg97=-114;	reg signed [w5-1:0] kh97=-69;	reg signed [w5-1:0] ki97=156;
reg signed [w5-1:0] ka98=-110;	reg signed [w5-1:0] kb98=-57;	reg signed [w5-1:0] kc98=-8;	reg signed [w5-1:0] kd98=108;	reg signed [w5-1:0] ke98=-142;	reg signed [w5-1:0] kf98=43;	reg signed [w5-1:0] kg98=-37;	reg signed [w5-1:0] kh98=75;	reg signed [w5-1:0] ki98=132;
reg signed [w5-1:0] ka99=-3;	reg signed [w5-1:0] kb99=157;	reg signed [w5-1:0] kc99=-54;	reg signed [w5-1:0] kd99=-138;	reg signed [w5-1:0] ke99=-114;	reg signed [w5-1:0] kf99=-113;	reg signed [w5-1:0] kg99=4;	reg signed [w5-1:0] kh99=-69;	reg signed [w5-1:0] ki99=31;
reg signed [w5-1:0] ka100=142;	reg signed [w5-1:0] kb100=76;	reg signed [w5-1:0] kc100=93;	reg signed [w5-1:0] kd100=137;	reg signed [w5-1:0] ke100=-98;	reg signed [w5-1:0] kf100=105;	reg signed [w5-1:0] kg100=89;	reg signed [w5-1:0] kh100=-87;	reg signed [w5-1:0] ki100=92;
reg signed [w5-1:0] ka101=77;	reg signed [w5-1:0] kb101=139;	reg signed [w5-1:0] kc101=23;	reg signed [w5-1:0] kd101=-141;	reg signed [w5-1:0] ke101=50;	reg signed [w5-1:0] kf101=178;	reg signed [w5-1:0] kg101=112;	reg signed [w5-1:0] kh101=-102;	reg signed [w5-1:0] ki101=129;
reg signed [w5-1:0] ka102=128;	reg signed [w5-1:0] kb102=-113;	reg signed [w5-1:0] kc102=-8;	reg signed [w5-1:0] kd102=-146;	reg signed [w5-1:0] ke102=-180;	reg signed [w5-1:0] kf102=-35;	reg signed [w5-1:0] kg102=70;	reg signed [w5-1:0] kh102=-175;	reg signed [w5-1:0] ki102=-19;
reg signed [w5-1:0] ka103=153;	reg signed [w5-1:0] kb103=8;	reg signed [w5-1:0] kc103=127;	reg signed [w5-1:0] kd103=94;	reg signed [w5-1:0] ke103=-50;	reg signed [w5-1:0] kf103=-137;	reg signed [w5-1:0] kg103=79;	reg signed [w5-1:0] kh103=-79;	reg signed [w5-1:0] ki103=109;
reg signed [w5-1:0] ka104=58;	reg signed [w5-1:0] kb104=-129;	reg signed [w5-1:0] kc104=190;	reg signed [w5-1:0] kd104=-46;	reg signed [w5-1:0] ke104=-95;	reg signed [w5-1:0] kf104=152;	reg signed [w5-1:0] kg104=45;	reg signed [w5-1:0] kh104=212;	reg signed [w5-1:0] ki104=150;
reg signed [w5-1:0] ka105=110;	reg signed [w5-1:0] kb105=-62;	reg signed [w5-1:0] kc105=-175;	reg signed [w5-1:0] kd105=92;	reg signed [w5-1:0] ke105=-11;	reg signed [w5-1:0] kf105=16;	reg signed [w5-1:0] kg105=2;	reg signed [w5-1:0] kh105=130;	reg signed [w5-1:0] ki105=-2;
reg signed [w5-1:0] ka106=-203;	reg signed [w5-1:0] kb106=48;	reg signed [w5-1:0] kc106=-12;	reg signed [w5-1:0] kd106=-10;	reg signed [w5-1:0] ke106=194;	reg signed [w5-1:0] kf106=160;	reg signed [w5-1:0] kg106=79;	reg signed [w5-1:0] kh106=120;	reg signed [w5-1:0] ki106=190;
reg signed [w5-1:0] ka107=15;	reg signed [w5-1:0] kb107=-17;	reg signed [w5-1:0] kc107=-69;	reg signed [w5-1:0] kd107=-34;	reg signed [w5-1:0] ke107=-129;	reg signed [w5-1:0] kf107=-189;	reg signed [w5-1:0] kg107=35;	reg signed [w5-1:0] kh107=23;	reg signed [w5-1:0] ki107=106;
reg signed [w5-1:0] ka108=-126;	reg signed [w5-1:0] kb108=-40;	reg signed [w5-1:0] kc108=-30;	reg signed [w5-1:0] kd108=-60;	reg signed [w5-1:0] ke108=-74;	reg signed [w5-1:0] kf108=-123;	reg signed [w5-1:0] kg108=71;	reg signed [w5-1:0] kh108=-58;	reg signed [w5-1:0] ki108=56;
reg signed [w5-1:0] ka109=10;	reg signed [w5-1:0] kb109=17;	reg signed [w5-1:0] kc109=-24;	reg signed [w5-1:0] kd109=31;	reg signed [w5-1:0] ke109=-47;	reg signed [w5-1:0] kf109=-63;	reg signed [w5-1:0] kg109=-80;	reg signed [w5-1:0] kh109=-122;	reg signed [w5-1:0] ki109=-4;
reg signed [w5-1:0] ka110=79;	reg signed [w5-1:0] kb110=-33;	reg signed [w5-1:0] kc110=-48;	reg signed [w5-1:0] kd110=49;	reg signed [w5-1:0] ke110=115;	reg signed [w5-1:0] kf110=86;	reg signed [w5-1:0] kg110=108;	reg signed [w5-1:0] kh110=19;	reg signed [w5-1:0] ki110=90;
reg signed [w5-1:0] ka111=7;	reg signed [w5-1:0] kb111=-93;	reg signed [w5-1:0] kc111=203;	reg signed [w5-1:0] kd111=-71;	reg signed [w5-1:0] ke111=-47;	reg signed [w5-1:0] kf111=72;	reg signed [w5-1:0] kg111=-12;	reg signed [w5-1:0] kh111=-106;	reg signed [w5-1:0] ki111=164;
reg signed [w5-1:0] ka112=-18;	reg signed [w5-1:0] kb112=22;	reg signed [w5-1:0] kc112=-101;	reg signed [w5-1:0] kd112=88;	reg signed [w5-1:0] ke112=112;	reg signed [w5-1:0] kf112=87;	reg signed [w5-1:0] kg112=-3;	reg signed [w5-1:0] kh112=-33;	reg signed [w5-1:0] ki112=55;
reg signed [w5-1:0] ka113=-72;	reg signed [w5-1:0] kb113=-170;	reg signed [w5-1:0] kc113=-174;	reg signed [w5-1:0] kd113=-37;	reg signed [w5-1:0] ke113=-84;	reg signed [w5-1:0] kf113=-144;	reg signed [w5-1:0] kg113=-29;	reg signed [w5-1:0] kh113=126;	reg signed [w5-1:0] ki113=30;
reg signed [w5-1:0] ka114=-119;	reg signed [w5-1:0] kb114=120;	reg signed [w5-1:0] kc114=67;	reg signed [w5-1:0] kd114=13;	reg signed [w5-1:0] ke114=-45;	reg signed [w5-1:0] kf114=60;	reg signed [w5-1:0] kg114=-131;	reg signed [w5-1:0] kh114=-14;	reg signed [w5-1:0] ki114=5;
reg signed [w5-1:0] ka115=-68;	reg signed [w5-1:0] kb115=-41;	reg signed [w5-1:0] kc115=110;	reg signed [w5-1:0] kd115=-53;	reg signed [w5-1:0] ke115=161;	reg signed [w5-1:0] kf115=-7;	reg signed [w5-1:0] kg115=139;	reg signed [w5-1:0] kh115=-42;	reg signed [w5-1:0] ki115=-13;
reg signed [w5-1:0] ka116=28;	reg signed [w5-1:0] kb116=174;	reg signed [w5-1:0] kc116=177;	reg signed [w5-1:0] kd116=145;	reg signed [w5-1:0] ke116=98;	reg signed [w5-1:0] kf116=95;	reg signed [w5-1:0] kg116=-34;	reg signed [w5-1:0] kh116=-131;	reg signed [w5-1:0] ki116=-45;
reg signed [w5-1:0] ka117=-43;	reg signed [w5-1:0] kb117=57;	reg signed [w5-1:0] kc117=-25;	reg signed [w5-1:0] kd117=-13;	reg signed [w5-1:0] ke117=79;	reg signed [w5-1:0] kf117=157;	reg signed [w5-1:0] kg117=-53;	reg signed [w5-1:0] kh117=73;	reg signed [w5-1:0] ki117=-51;
reg signed [w5-1:0] ka118=119;	reg signed [w5-1:0] kb118=90;	reg signed [w5-1:0] kc118=56;	reg signed [w5-1:0] kd118=-123;	reg signed [w5-1:0] ke118=112;	reg signed [w5-1:0] kf118=84;	reg signed [w5-1:0] kg118=-43;	reg signed [w5-1:0] kh118=-42;	reg signed [w5-1:0] ki118=59;
reg signed [w5-1:0] ka119=-35;	reg signed [w5-1:0] kb119=15;	reg signed [w5-1:0] kc119=98;	reg signed [w5-1:0] kd119=12;	reg signed [w5-1:0] ke119=3;	reg signed [w5-1:0] kf119=-112;	reg signed [w5-1:0] kg119=136;	reg signed [w5-1:0] kh119=129;	reg signed [w5-1:0] ki119=-30;
reg signed [w5-1:0] ka120=-172;	reg signed [w5-1:0] kb120=-152;	reg signed [w5-1:0] kc120=-84;	reg signed [w5-1:0] kd120=5;	reg signed [w5-1:0] ke120=101;	reg signed [w5-1:0] kf120=-76;	reg signed [w5-1:0] kg120=190;	reg signed [w5-1:0] kh120=-132;	reg signed [w5-1:0] ki120=-67;
reg signed [w5-1:0] ka121=14;	reg signed [w5-1:0] kb121=67;	reg signed [w5-1:0] kc121=0;	reg signed [w5-1:0] kd121=-71;	reg signed [w5-1:0] ke121=-56;	reg signed [w5-1:0] kf121=-9;	reg signed [w5-1:0] kg121=-125;	reg signed [w5-1:0] kh121=-22;	reg signed [w5-1:0] ki121=-46;
reg signed [w5-1:0] ka122=-49;	reg signed [w5-1:0] kb122=-118;	reg signed [w5-1:0] kc122=54;	reg signed [w5-1:0] kd122=-38;	reg signed [w5-1:0] ke122=-97;	reg signed [w5-1:0] kf122=-16;	reg signed [w5-1:0] kg122=-50;	reg signed [w5-1:0] kh122=-129;	reg signed [w5-1:0] ki122=82;
reg signed [w5-1:0] ka123=101;	reg signed [w5-1:0] kb123=-76;	reg signed [w5-1:0] kc123=102;	reg signed [w5-1:0] kd123=-96;	reg signed [w5-1:0] ke123=-23;	reg signed [w5-1:0] kf123=-32;	reg signed [w5-1:0] kg123=-102;	reg signed [w5-1:0] kh123=64;	reg signed [w5-1:0] ki123=-170;
reg signed [w5-1:0] ka124=99;	reg signed [w5-1:0] kb124=-14;	reg signed [w5-1:0] kc124=30;	reg signed [w5-1:0] kd124=-94;	reg signed [w5-1:0] ke124=-139;	reg signed [w5-1:0] kf124=45;	reg signed [w5-1:0] kg124=-14;	reg signed [w5-1:0] kh124=-41;	reg signed [w5-1:0] ki124=87;
reg signed [w5-1:0] ka125=304;	reg signed [w5-1:0] kb125=65;	reg signed [w5-1:0] kc125=-43;	reg signed [w5-1:0] kd125=-112;	reg signed [w5-1:0] ke125=83;	reg signed [w5-1:0] kf125=-84;	reg signed [w5-1:0] kg125=25;	reg signed [w5-1:0] kh125=-88;	reg signed [w5-1:0] ki125=-99;
reg signed [w5-1:0] ka126=-13;	reg signed [w5-1:0] kb126=105;	reg signed [w5-1:0] kc126=-165;	reg signed [w5-1:0] kd126=-137;	reg signed [w5-1:0] ke126=-58;	reg signed [w5-1:0] kf126=46;	reg signed [w5-1:0] kg126=24;	reg signed [w5-1:0] kh126=25;	reg signed [w5-1:0] ki126=51;
reg signed [w5-1:0] ka127=-47;	reg signed [w5-1:0] kb127=-3;	reg signed [w5-1:0] kc127=-83;	reg signed [w5-1:0] kd127=141;	reg signed [w5-1:0] ke127=-69;	reg signed [w5-1:0] kf127=16;	reg signed [w5-1:0] kg127=-22;	reg signed [w5-1:0] kh127=128;	reg signed [w5-1:0] ki127=56;
reg signed [w5-1:0] ka128=185;	reg signed [w5-1:0] kb128=161;	reg signed [w5-1:0] kc128=-127;	reg signed [w5-1:0] kd128=146;	reg signed [w5-1:0] ke128=48;	reg signed [w5-1:0] kf128=-50;	reg signed [w5-1:0] kg128=-146;	reg signed [w5-1:0] kh128=-153;	reg signed [w5-1:0] ki128=-55;
reg signed [w5-1:0] ka129=75;	reg signed [w5-1:0] kb129=191;	reg signed [w5-1:0] kc129=119;	reg signed [w5-1:0] kd129=141;	reg signed [w5-1:0] ke129=106;	reg signed [w5-1:0] kf129=102;	reg signed [w5-1:0] kg129=74;	reg signed [w5-1:0] kh129=4;	reg signed [w5-1:0] ki129=-136;
reg signed [w5-1:0] ka130=81;	reg signed [w5-1:0] kb130=34;	reg signed [w5-1:0] kc130=38;	reg signed [w5-1:0] kd130=-14;	reg signed [w5-1:0] ke130=-206;	reg signed [w5-1:0] kf130=-46;	reg signed [w5-1:0] kg130=-73;	reg signed [w5-1:0] kh130=-118;	reg signed [w5-1:0] ki130=41;
reg signed [w5-1:0] ka131=133;	reg signed [w5-1:0] kb131=86;	reg signed [w5-1:0] kc131=40;	reg signed [w5-1:0] kd131=-47;	reg signed [w5-1:0] ke131=-17;	reg signed [w5-1:0] kf131=92;	reg signed [w5-1:0] kg131=71;	reg signed [w5-1:0] kh131=39;	reg signed [w5-1:0] ki131=55;
reg signed [w5-1:0] ka132=-41;	reg signed [w5-1:0] kb132=195;	reg signed [w5-1:0] kc132=53;	reg signed [w5-1:0] kd132=-55;	reg signed [w5-1:0] ke132=178;	reg signed [w5-1:0] kf132=-98;	reg signed [w5-1:0] kg132=80;	reg signed [w5-1:0] kh132=177;	reg signed [w5-1:0] ki132=44;
reg signed [w5-1:0] ka133=-104;	reg signed [w5-1:0] kb133=-131;	reg signed [w5-1:0] kc133=-56;	reg signed [w5-1:0] kd133=124;	reg signed [w5-1:0] ke133=7;	reg signed [w5-1:0] kf133=20;	reg signed [w5-1:0] kg133=147;	reg signed [w5-1:0] kh133=113;	reg signed [w5-1:0] ki133=-139;
reg signed [w5-1:0] ka134=-30;	reg signed [w5-1:0] kb134=-189;	reg signed [w5-1:0] kc134=33;	reg signed [w5-1:0] kd134=-41;	reg signed [w5-1:0] ke134=64;	reg signed [w5-1:0] kf134=125;	reg signed [w5-1:0] kg134=46;	reg signed [w5-1:0] kh134=-87;	reg signed [w5-1:0] ki134=178;
reg signed [w5-1:0] ka135=148;	reg signed [w5-1:0] kb135=-127;	reg signed [w5-1:0] kc135=-196;	reg signed [w5-1:0] kd135=-98;	reg signed [w5-1:0] ke135=69;	reg signed [w5-1:0] kf135=13;	reg signed [w5-1:0] kg135=31;	reg signed [w5-1:0] kh135=40;	reg signed [w5-1:0] ki135=190;
reg signed [w5-1:0] ka136=109;	reg signed [w5-1:0] kb136=-48;	reg signed [w5-1:0] kc136=-162;	reg signed [w5-1:0] kd136=76;	reg signed [w5-1:0] ke136=-116;	reg signed [w5-1:0] kf136=-144;	reg signed [w5-1:0] kg136=94;	reg signed [w5-1:0] kh136=-32;	reg signed [w5-1:0] ki136=-77;

reg signed [w7-1:0] delta9=1265;	reg signed [w7-1:0] mu9=-126;	reg signed [w7-1:0] beta9=-11039;
reg signed [w7-1:0] delta10=961;	reg signed [w7-1:0] mu10=962;	reg signed [w7-1:0] beta10=-15035;
reg signed [w7-1:0] delta11=1219;	reg signed [w7-1:0] mu11=233;	reg signed [w7-1:0] beta11=-25538;
reg signed [w7-1:0] delta12=1592;	reg signed [w7-1:0] mu12=-104;	reg signed [w7-1:0] beta12=-1310;
reg signed [w7-1:0] delta13=1225;	reg signed [w7-1:0] mu13=277;	reg signed [w7-1:0] beta13=-20787;
reg signed [w7-1:0] delta14=1997;	reg signed [w7-1:0] mu14=409;	reg signed [w7-1:0] beta14=6421;
reg signed [w7-1:0] delta15=1181;	reg signed [w7-1:0] mu15=998;	reg signed [w7-1:0] beta15=21653;
reg signed [w7-1:0] delta16=1214;	reg signed [w7-1:0] mu16=186;	reg signed [w7-1:0] beta16=7653;
reg signed [w7-1:0] delta17=1291;	reg signed [w7-1:0] mu17=661;	reg signed [w7-1:0] beta17=12072;
reg signed [w7-1:0] delta18=1546;	reg signed [w7-1:0] mu18=20;	reg signed [w7-1:0] beta18=-32843;
reg signed [w7-1:0] delta19=1215;	reg signed [w7-1:0] mu19=-596;	reg signed [w7-1:0] beta19=-19119;
reg signed [w7-1:0] delta20=1490;	reg signed [w7-1:0] mu20=302;	reg signed [w7-1:0] beta20=-4934;
reg signed [w7-1:0] delta21=1249;	reg signed [w7-1:0] mu21=199;	reg signed [w7-1:0] beta21=13226;
reg signed [w7-1:0] delta22=1160;	reg signed [w7-1:0] mu22=275;	reg signed [w7-1:0] beta22=-27932;
reg signed [w7-1:0] delta23=1605;	reg signed [w7-1:0] mu23=-391;	reg signed [w7-1:0] beta23=-82773;
reg signed [w7-1:0] delta24=1159;	reg signed [w7-1:0] mu24=603;	reg signed [w7-1:0] beta24=4530;


reg signed [w10-1:0] ka137=85;	reg signed [w10-1:0] kb137=20;	reg signed [w10-1:0] kc137=35;	reg signed [w10-1:0] kd137=98;	reg signed [w10-1:0] ke137=101;	reg signed [w10-1:0] kf137=-124;	reg signed [w10-1:0] kg137=-55;	reg signed [w10-1:0] kh137=-79;	reg signed [w10-1:0] ki137=97;
reg signed [w10-1:0] ka138=-25;	reg signed [w10-1:0] kb138=16;	reg signed [w10-1:0] kc138=-16;	reg signed [w10-1:0] kd138=102;	reg signed [w10-1:0] ke138=-130;	reg signed [w10-1:0] kf138=-89;	reg signed [w10-1:0] kg138=65;	reg signed [w10-1:0] kh138=-68;	reg signed [w10-1:0] ki138=47;
reg signed [w10-1:0] ka139=114;	reg signed [w10-1:0] kb139=-6;	reg signed [w10-1:0] kc139=-132;	reg signed [w10-1:0] kd139=-27;	reg signed [w10-1:0] ke139=55;	reg signed [w10-1:0] kf139=-42;	reg signed [w10-1:0] kg139=-100;	reg signed [w10-1:0] kh139=31;	reg signed [w10-1:0] ki139=52;
reg signed [w10-1:0] ka140=-13;	reg signed [w10-1:0] kb140=98;	reg signed [w10-1:0] kc140=-27;	reg signed [w10-1:0] kd140=109;	reg signed [w10-1:0] ke140=36;	reg signed [w10-1:0] kf140=110;	reg signed [w10-1:0] kg140=-72;	reg signed [w10-1:0] kh140=-84;	reg signed [w10-1:0] ki140=-4;
reg signed [w10-1:0] ka141=8;	reg signed [w10-1:0] kb141=-42;	reg signed [w10-1:0] kc141=23;	reg signed [w10-1:0] kd141=-31;	reg signed [w10-1:0] ke141=5;	reg signed [w10-1:0] kf141=143;	reg signed [w10-1:0] kg141=-54;	reg signed [w10-1:0] kh141=109;	reg signed [w10-1:0] ki141=-19;
reg signed [w10-1:0] ka142=74;	reg signed [w10-1:0] kb142=48;	reg signed [w10-1:0] kc142=68;	reg signed [w10-1:0] kd142=14;	reg signed [w10-1:0] ke142=-86;	reg signed [w10-1:0] kf142=-79;	reg signed [w10-1:0] kg142=43;	reg signed [w10-1:0] kh142=-65;	reg signed [w10-1:0] ki142=-80;
reg signed [w10-1:0] ka143=-40;	reg signed [w10-1:0] kb143=45;	reg signed [w10-1:0] kc143=-11;	reg signed [w10-1:0] kd143=150;	reg signed [w10-1:0] ke143=-14;	reg signed [w10-1:0] kf143=77;	reg signed [w10-1:0] kg143=-15;	reg signed [w10-1:0] kh143=110;	reg signed [w10-1:0] ki143=-102;
reg signed [w10-1:0] ka144=-56;	reg signed [w10-1:0] kb144=-153;	reg signed [w10-1:0] kc144=-67;	reg signed [w10-1:0] kd144=75;	reg signed [w10-1:0] ke144=-17;	reg signed [w10-1:0] kf144=-75;	reg signed [w10-1:0] kg144=-67;	reg signed [w10-1:0] kh144=-86;	reg signed [w10-1:0] ki144=-49;
reg signed [w10-1:0] ka145=85;	reg signed [w10-1:0] kb145=139;	reg signed [w10-1:0] kc145=46;	reg signed [w10-1:0] kd145=35;	reg signed [w10-1:0] ke145=-127;	reg signed [w10-1:0] kf145=76;	reg signed [w10-1:0] kg145=-35;	reg signed [w10-1:0] kh145=-103;	reg signed [w10-1:0] ki145=-24;
reg signed [w10-1:0] ka146=87;	reg signed [w10-1:0] kb146=157;	reg signed [w10-1:0] kc146=182;	reg signed [w10-1:0] kd146=13;	reg signed [w10-1:0] ke146=-5;	reg signed [w10-1:0] kf146=127;	reg signed [w10-1:0] kg146=-121;	reg signed [w10-1:0] kh146=14;	reg signed [w10-1:0] ki146=56;
reg signed [w10-1:0] ka147=-71;	reg signed [w10-1:0] kb147=-59;	reg signed [w10-1:0] kc147=-36;	reg signed [w10-1:0] kd147=-16;	reg signed [w10-1:0] ke147=-25;	reg signed [w10-1:0] kf147=-106;	reg signed [w10-1:0] kg147=35;	reg signed [w10-1:0] kh147=35;	reg signed [w10-1:0] ki147=9;
reg signed [w10-1:0] ka148=19;	reg signed [w10-1:0] kb148=60;	reg signed [w10-1:0] kc148=122;	reg signed [w10-1:0] kd148=50;	reg signed [w10-1:0] ke148=34;	reg signed [w10-1:0] kf148=158;	reg signed [w10-1:0] kg148=102;	reg signed [w10-1:0] kh148=21;	reg signed [w10-1:0] ki148=145;
reg signed [w10-1:0] ka149=-59;	reg signed [w10-1:0] kb149=-13;	reg signed [w10-1:0] kc149=6;	reg signed [w10-1:0] kd149=117;	reg signed [w10-1:0] ke149=1;	reg signed [w10-1:0] kf149=-55;	reg signed [w10-1:0] kg149=85;	reg signed [w10-1:0] kh149=-30;	reg signed [w10-1:0] ki149=87;
reg signed [w10-1:0] ka150=-63;	reg signed [w10-1:0] kb150=31;	reg signed [w10-1:0] kc150=62;	reg signed [w10-1:0] kd150=92;	reg signed [w10-1:0] ke150=71;	reg signed [w10-1:0] kf150=-118;	reg signed [w10-1:0] kg150=39;	reg signed [w10-1:0] kh150=70;	reg signed [w10-1:0] ki150=98;
reg signed [w10-1:0] ka151=15;	reg signed [w10-1:0] kb151=101;	reg signed [w10-1:0] kc151=40;	reg signed [w10-1:0] kd151=-51;	reg signed [w10-1:0] ke151=37;	reg signed [w10-1:0] kf151=-95;	reg signed [w10-1:0] kg151=34;	reg signed [w10-1:0] kh151=-45;	reg signed [w10-1:0] ki151=-51;
reg signed [w10-1:0] ka152=-119;	reg signed [w10-1:0] kb152=-136;	reg signed [w10-1:0] kc152=-146;	reg signed [w10-1:0] kd152=70;	reg signed [w10-1:0] ke152=-54;	reg signed [w10-1:0] kf152=-9;	reg signed [w10-1:0] kg152=-80;	reg signed [w10-1:0] kh152=72;	reg signed [w10-1:0] ki152=-16;
reg signed [w10-1:0] ka153=-72;	reg signed [w10-1:0] kb153=22;	reg signed [w10-1:0] kc153=-56;	reg signed [w10-1:0] kd153=-24;	reg signed [w10-1:0] ke153=65;	reg signed [w10-1:0] kf153=-54;	reg signed [w10-1:0] kg153=-107;	reg signed [w10-1:0] kh153=11;	reg signed [w10-1:0] ki153=-40;
reg signed [w10-1:0] ka154=22;	reg signed [w10-1:0] kb154=-70;	reg signed [w10-1:0] kc154=25;	reg signed [w10-1:0] kd154=55;	reg signed [w10-1:0] ke154=-112;	reg signed [w10-1:0] kf154=-132;	reg signed [w10-1:0] kg154=38;	reg signed [w10-1:0] kh154=-47;	reg signed [w10-1:0] ki154=-1;
reg signed [w10-1:0] ka155=122;	reg signed [w10-1:0] kb155=47;	reg signed [w10-1:0] kc155=45;	reg signed [w10-1:0] kd155=72;	reg signed [w10-1:0] ke155=60;	reg signed [w10-1:0] kf155=-73;	reg signed [w10-1:0] kg155=-26;	reg signed [w10-1:0] kh155=73;	reg signed [w10-1:0] ki155=55;
reg signed [w10-1:0] ka156=-29;	reg signed [w10-1:0] kb156=-87;	reg signed [w10-1:0] kc156=27;	reg signed [w10-1:0] kd156=61;	reg signed [w10-1:0] ke156=89;	reg signed [w10-1:0] kf156=43;	reg signed [w10-1:0] kg156=-57;	reg signed [w10-1:0] kh156=28;	reg signed [w10-1:0] ki156=4;
reg signed [w10-1:0] ka157=-46;	reg signed [w10-1:0] kb157=-12;	reg signed [w10-1:0] kc157=-113;	reg signed [w10-1:0] kd157=21;	reg signed [w10-1:0] ke157=-24;	reg signed [w10-1:0] kf157=125;	reg signed [w10-1:0] kg157=-117;	reg signed [w10-1:0] kh157=93;	reg signed [w10-1:0] ki157=88;
reg signed [w10-1:0] ka158=-60;	reg signed [w10-1:0] kb158=-10;	reg signed [w10-1:0] kc158=-141;	reg signed [w10-1:0] kd158=50;	reg signed [w10-1:0] ke158=-20;	reg signed [w10-1:0] kf158=-47;	reg signed [w10-1:0] kg158=4;	reg signed [w10-1:0] kh158=-72;	reg signed [w10-1:0] ki158=-121;
reg signed [w10-1:0] ka159=41;	reg signed [w10-1:0] kb159=88;	reg signed [w10-1:0] kc159=-29;	reg signed [w10-1:0] kd159=46;	reg signed [w10-1:0] ke159=114;	reg signed [w10-1:0] kf159=-8;	reg signed [w10-1:0] kg159=-130;	reg signed [w10-1:0] kh159=3;	reg signed [w10-1:0] ki159=-107;
reg signed [w10-1:0] ka160=-4;	reg signed [w10-1:0] kb160=-118;	reg signed [w10-1:0] kc160=-32;	reg signed [w10-1:0] kd160=-98;	reg signed [w10-1:0] ke160=-32;	reg signed [w10-1:0] kf160=145;	reg signed [w10-1:0] kg160=49;	reg signed [w10-1:0] kh160=-14;	reg signed [w10-1:0] ki160=202;
reg signed [w10-1:0] ka161=-99;	reg signed [w10-1:0] kb161=-20;	reg signed [w10-1:0] kc161=113;	reg signed [w10-1:0] kd161=91;	reg signed [w10-1:0] ke161=108;	reg signed [w10-1:0] kf161=-66;	reg signed [w10-1:0] kg161=12;	reg signed [w10-1:0] kh161=85;	reg signed [w10-1:0] ki161=63;
reg signed [w10-1:0] ka162=-11;	reg signed [w10-1:0] kb162=-39;	reg signed [w10-1:0] kc162=4;	reg signed [w10-1:0] kd162=-6;	reg signed [w10-1:0] ke162=-27;	reg signed [w10-1:0] kf162=31;	reg signed [w10-1:0] kg162=92;	reg signed [w10-1:0] kh162=-116;	reg signed [w10-1:0] ki162=-88;
reg signed [w10-1:0] ka163=-31;	reg signed [w10-1:0] kb163=50;	reg signed [w10-1:0] kc163=51;	reg signed [w10-1:0] kd163=28;	reg signed [w10-1:0] ke163=-89;	reg signed [w10-1:0] kf163=12;	reg signed [w10-1:0] kg163=87;	reg signed [w10-1:0] kh163=-22;	reg signed [w10-1:0] ki163=-81;
reg signed [w10-1:0] ka164=-56;	reg signed [w10-1:0] kb164=106;	reg signed [w10-1:0] kc164=62;	reg signed [w10-1:0] kd164=94;	reg signed [w10-1:0] ke164=-9;	reg signed [w10-1:0] kf164=-47;	reg signed [w10-1:0] kg164=145;	reg signed [w10-1:0] kh164=-15;	reg signed [w10-1:0] ki164=-58;
reg signed [w10-1:0] ka165=87;	reg signed [w10-1:0] kb165=61;	reg signed [w10-1:0] kc165=-92;	reg signed [w10-1:0] kd165=73;	reg signed [w10-1:0] ke165=-29;	reg signed [w10-1:0] kf165=-127;	reg signed [w10-1:0] kg165=-72;	reg signed [w10-1:0] kh165=-148;	reg signed [w10-1:0] ki165=23;
reg signed [w10-1:0] ka166=15;	reg signed [w10-1:0] kb166=25;	reg signed [w10-1:0] kc166=-21;	reg signed [w10-1:0] kd166=-60;	reg signed [w10-1:0] ke166=-36;	reg signed [w10-1:0] kf166=85;	reg signed [w10-1:0] kg166=22;	reg signed [w10-1:0] kh166=-75;	reg signed [w10-1:0] ki166=69;
reg signed [w10-1:0] ka167=42;	reg signed [w10-1:0] kb167=-40;	reg signed [w10-1:0] kc167=-56;	reg signed [w10-1:0] kd167=17;	reg signed [w10-1:0] ke167=-126;	reg signed [w10-1:0] kf167=-63;	reg signed [w10-1:0] kg167=10;	reg signed [w10-1:0] kh167=42;	reg signed [w10-1:0] ki167=-63;
reg signed [w10-1:0] ka168=11;	reg signed [w10-1:0] kb168=-123;	reg signed [w10-1:0] kc168=4;	reg signed [w10-1:0] kd168=-118;	reg signed [w10-1:0] ke168=-4;	reg signed [w10-1:0] kf168=140;	reg signed [w10-1:0] kg168=-85;	reg signed [w10-1:0] kh168=-47;	reg signed [w10-1:0] ki168=-39;
reg signed [w10-1:0] ka169=-62;	reg signed [w10-1:0] kb169=-28;	reg signed [w10-1:0] kc169=43;	reg signed [w10-1:0] kd169=-75;	reg signed [w10-1:0] ke169=-104;	reg signed [w10-1:0] kf169=-10;	reg signed [w10-1:0] kg169=-22;	reg signed [w10-1:0] kh169=-55;	reg signed [w10-1:0] ki169=-23;
reg signed [w10-1:0] ka170=77;	reg signed [w10-1:0] kb170=27;	reg signed [w10-1:0] kc170=35;	reg signed [w10-1:0] kd170=45;	reg signed [w10-1:0] ke170=112;	reg signed [w10-1:0] kf170=50;	reg signed [w10-1:0] kg170=-67;	reg signed [w10-1:0] kh170=6;	reg signed [w10-1:0] ki170=-80;
reg signed [w10-1:0] ka171=30;	reg signed [w10-1:0] kb171=23;	reg signed [w10-1:0] kc171=81;	reg signed [w10-1:0] kd171=-72;	reg signed [w10-1:0] ke171=-38;	reg signed [w10-1:0] kf171=-15;	reg signed [w10-1:0] kg171=38;	reg signed [w10-1:0] kh171=-41;	reg signed [w10-1:0] ki171=-30;
reg signed [w10-1:0] ka172=37;	reg signed [w10-1:0] kb172=-90;	reg signed [w10-1:0] kc172=-40;	reg signed [w10-1:0] kd172=29;	reg signed [w10-1:0] ke172=20;	reg signed [w10-1:0] kf172=31;	reg signed [w10-1:0] kg172=9;	reg signed [w10-1:0] kh172=82;	reg signed [w10-1:0] ki172=112;
reg signed [w10-1:0] ka173=38;	reg signed [w10-1:0] kb173=-79;	reg signed [w10-1:0] kc173=3;	reg signed [w10-1:0] kd173=30;	reg signed [w10-1:0] ke173=-96;	reg signed [w10-1:0] kf173=83;	reg signed [w10-1:0] kg173=19;	reg signed [w10-1:0] kh173=-64;	reg signed [w10-1:0] ki173=-2;
reg signed [w10-1:0] ka174=69;	reg signed [w10-1:0] kb174=114;	reg signed [w10-1:0] kc174=81;	reg signed [w10-1:0] kd174=-107;	reg signed [w10-1:0] ke174=-117;	reg signed [w10-1:0] kf174=25;	reg signed [w10-1:0] kg174=-48;	reg signed [w10-1:0] kh174=2;	reg signed [w10-1:0] ki174=50;
reg signed [w10-1:0] ka175=29;	reg signed [w10-1:0] kb175=100;	reg signed [w10-1:0] kc175=107;	reg signed [w10-1:0] kd175=89;	reg signed [w10-1:0] ke175=78;	reg signed [w10-1:0] kf175=151;	reg signed [w10-1:0] kg175=50;	reg signed [w10-1:0] kh175=97;	reg signed [w10-1:0] ki175=84;
reg signed [w10-1:0] ka176=-13;	reg signed [w10-1:0] kb176=-95;	reg signed [w10-1:0] kc176=7;	reg signed [w10-1:0] kd176=-109;	reg signed [w10-1:0] ke176=-120;	reg signed [w10-1:0] kf176=-70;	reg signed [w10-1:0] kg176=106;	reg signed [w10-1:0] kh176=53;	reg signed [w10-1:0] ki176=-34;
reg signed [w10-1:0] ka177=119;	reg signed [w10-1:0] kb177=46;	reg signed [w10-1:0] kc177=-72;	reg signed [w10-1:0] kd177=65;	reg signed [w10-1:0] ke177=-51;	reg signed [w10-1:0] kf177=-18;	reg signed [w10-1:0] kg177=2;	reg signed [w10-1:0] kh177=-15;	reg signed [w10-1:0] ki177=157;
reg signed [w10-1:0] ka178=16;	reg signed [w10-1:0] kb178=-76;	reg signed [w10-1:0] kc178=-6;	reg signed [w10-1:0] kd178=79;	reg signed [w10-1:0] ke178=58;	reg signed [w10-1:0] kf178=-122;	reg signed [w10-1:0] kg178=-26;	reg signed [w10-1:0] kh178=176;	reg signed [w10-1:0] ki178=197;
reg signed [w10-1:0] ka179=113;	reg signed [w10-1:0] kb179=-21;	reg signed [w10-1:0] kc179=-57;	reg signed [w10-1:0] kd179=-68;	reg signed [w10-1:0] ke179=-79;	reg signed [w10-1:0] kf179=-16;	reg signed [w10-1:0] kg179=103;	reg signed [w10-1:0] kh179=-85;	reg signed [w10-1:0] ki179=-94;
reg signed [w10-1:0] ka180=97;	reg signed [w10-1:0] kb180=6;	reg signed [w10-1:0] kc180=52;	reg signed [w10-1:0] kd180=-47;	reg signed [w10-1:0] ke180=136;	reg signed [w10-1:0] kf180=81;	reg signed [w10-1:0] kg180=-27;	reg signed [w10-1:0] kh180=-48;	reg signed [w10-1:0] ki180=16;
reg signed [w10-1:0] ka181=-22;	reg signed [w10-1:0] kb181=64;	reg signed [w10-1:0] kc181=66;	reg signed [w10-1:0] kd181=-83;	reg signed [w10-1:0] ke181=21;	reg signed [w10-1:0] kf181=-29;	reg signed [w10-1:0] kg181=-50;	reg signed [w10-1:0] kh181=-111;	reg signed [w10-1:0] ki181=50;
reg signed [w10-1:0] ka182=20;	reg signed [w10-1:0] kb182=57;	reg signed [w10-1:0] kc182=113;	reg signed [w10-1:0] kd182=-124;	reg signed [w10-1:0] ke182=-74;	reg signed [w10-1:0] kf182=-12;	reg signed [w10-1:0] kg182=-131;	reg signed [w10-1:0] kh182=-55;	reg signed [w10-1:0] ki182=-75;
reg signed [w10-1:0] ka183=34;	reg signed [w10-1:0] kb183=-1;	reg signed [w10-1:0] kc183=40;	reg signed [w10-1:0] kd183=-34;	reg signed [w10-1:0] ke183=9;	reg signed [w10-1:0] kf183=-148;	reg signed [w10-1:0] kg183=-76;	reg signed [w10-1:0] kh183=100;	reg signed [w10-1:0] ki183=-131;
reg signed [w10-1:0] ka184=-50;	reg signed [w10-1:0] kb184=-98;	reg signed [w10-1:0] kc184=-20;	reg signed [w10-1:0] kd184=87;	reg signed [w10-1:0] ke184=94;	reg signed [w10-1:0] kf184=-64;	reg signed [w10-1:0] kg184=63;	reg signed [w10-1:0] kh184=-65;	reg signed [w10-1:0] ki184=-14;
reg signed [w10-1:0] ka185=-80;	reg signed [w10-1:0] kb185=-73;	reg signed [w10-1:0] kc185=146;	reg signed [w10-1:0] kd185=13;	reg signed [w10-1:0] ke185=133;	reg signed [w10-1:0] kf185=45;	reg signed [w10-1:0] kg185=-31;	reg signed [w10-1:0] kh185=-101;	reg signed [w10-1:0] ki185=69;
reg signed [w10-1:0] ka186=102;	reg signed [w10-1:0] kb186=-14;	reg signed [w10-1:0] kc186=8;	reg signed [w10-1:0] kd186=-104;	reg signed [w10-1:0] ke186=-93;	reg signed [w10-1:0] kf186=101;	reg signed [w10-1:0] kg186=41;	reg signed [w10-1:0] kh186=33;	reg signed [w10-1:0] ki186=84;
reg signed [w10-1:0] ka187=-65;	reg signed [w10-1:0] kb187=72;	reg signed [w10-1:0] kc187=8;	reg signed [w10-1:0] kd187=58;	reg signed [w10-1:0] ke187=85;	reg signed [w10-1:0] kf187=118;	reg signed [w10-1:0] kg187=63;	reg signed [w10-1:0] kh187=2;	reg signed [w10-1:0] ki187=146;
reg signed [w10-1:0] ka188=41;	reg signed [w10-1:0] kb188=61;	reg signed [w10-1:0] kc188=-48;	reg signed [w10-1:0] kd188=4;	reg signed [w10-1:0] ke188=-54;	reg signed [w10-1:0] kf188=68;	reg signed [w10-1:0] kg188=59;	reg signed [w10-1:0] kh188=-22;	reg signed [w10-1:0] ki188=-97;
reg signed [w10-1:0] ka189=-41;	reg signed [w10-1:0] kb189=-33;	reg signed [w10-1:0] kc189=-15;	reg signed [w10-1:0] kd189=24;	reg signed [w10-1:0] ke189=-45;	reg signed [w10-1:0] kf189=-64;	reg signed [w10-1:0] kg189=30;	reg signed [w10-1:0] kh189=-6;	reg signed [w10-1:0] ki189=-80;
reg signed [w10-1:0] ka190=1;	reg signed [w10-1:0] kb190=-23;	reg signed [w10-1:0] kc190=-116;	reg signed [w10-1:0] kd190=37;	reg signed [w10-1:0] ke190=-69;	reg signed [w10-1:0] kf190=-73;	reg signed [w10-1:0] kg190=46;	reg signed [w10-1:0] kh190=-93;	reg signed [w10-1:0] ki190=-24;
reg signed [w10-1:0] ka191=-20;	reg signed [w10-1:0] kb191=27;	reg signed [w10-1:0] kc191=-84;	reg signed [w10-1:0] kd191=-14;	reg signed [w10-1:0] ke191=-71;	reg signed [w10-1:0] kf191=-32;	reg signed [w10-1:0] kg191=49;	reg signed [w10-1:0] kh191=28;	reg signed [w10-1:0] ki191=-26;
reg signed [w10-1:0] ka192=18;	reg signed [w10-1:0] kb192=-56;	reg signed [w10-1:0] kc192=-72;	reg signed [w10-1:0] kd192=-91;	reg signed [w10-1:0] ke192=-71;	reg signed [w10-1:0] kf192=-44;	reg signed [w10-1:0] kg192=141;	reg signed [w10-1:0] kh192=-106;	reg signed [w10-1:0] ki192=-24;
reg signed [w10-1:0] ka193=80;	reg signed [w10-1:0] kb193=46;	reg signed [w10-1:0] kc193=1;	reg signed [w10-1:0] kd193=-39;	reg signed [w10-1:0] ke193=53;	reg signed [w10-1:0] kf193=69;	reg signed [w10-1:0] kg193=-102;	reg signed [w10-1:0] kh193=33;	reg signed [w10-1:0] ki193=-36;
reg signed [w10-1:0] ka194=-60;	reg signed [w10-1:0] kb194=28;	reg signed [w10-1:0] kc194=-51;	reg signed [w10-1:0] kd194=3;	reg signed [w10-1:0] ke194=38;	reg signed [w10-1:0] kf194=-44;	reg signed [w10-1:0] kg194=-37;	reg signed [w10-1:0] kh194=-112;	reg signed [w10-1:0] ki194=135;
reg signed [w10-1:0] ka195=70;	reg signed [w10-1:0] kb195=68;	reg signed [w10-1:0] kc195=73;	reg signed [w10-1:0] kd195=-40;	reg signed [w10-1:0] ke195=18;	reg signed [w10-1:0] kf195=12;	reg signed [w10-1:0] kg195=48;	reg signed [w10-1:0] kh195=102;	reg signed [w10-1:0] ki195=-81;
reg signed [w10-1:0] ka196=120;	reg signed [w10-1:0] kb196=-17;	reg signed [w10-1:0] kc196=109;	reg signed [w10-1:0] kd196=-83;	reg signed [w10-1:0] ke196=71;	reg signed [w10-1:0] kf196=92;	reg signed [w10-1:0] kg196=-12;	reg signed [w10-1:0] kh196=88;	reg signed [w10-1:0] ki196=-105;
reg signed [w10-1:0] ka197=40;	reg signed [w10-1:0] kb197=15;	reg signed [w10-1:0] kc197=-28;	reg signed [w10-1:0] kd197=-24;	reg signed [w10-1:0] ke197=-11;	reg signed [w10-1:0] kf197=-133;	reg signed [w10-1:0] kg197=-75;	reg signed [w10-1:0] kh197=-58;	reg signed [w10-1:0] ki197=-94;
reg signed [w10-1:0] ka198=-51;	reg signed [w10-1:0] kb198=-110;	reg signed [w10-1:0] kc198=38;	reg signed [w10-1:0] kd198=26;	reg signed [w10-1:0] ke198=-147;	reg signed [w10-1:0] kf198=-85;	reg signed [w10-1:0] kg198=-42;	reg signed [w10-1:0] kh198=87;	reg signed [w10-1:0] ki198=97;
reg signed [w10-1:0] ka199=-50;	reg signed [w10-1:0] kb199=-55;	reg signed [w10-1:0] kc199=-96;	reg signed [w10-1:0] kd199=-100;	reg signed [w10-1:0] ke199=-118;	reg signed [w10-1:0] kf199=-50;	reg signed [w10-1:0] kg199=29;	reg signed [w10-1:0] kh199=-71;	reg signed [w10-1:0] ki199=-43;
reg signed [w10-1:0] ka200=-132;	reg signed [w10-1:0] kb200=-27;	reg signed [w10-1:0] kc200=-73;	reg signed [w10-1:0] kd200=-21;	reg signed [w10-1:0] ke200=125;	reg signed [w10-1:0] kf200=143;	reg signed [w10-1:0] kg200=46;	reg signed [w10-1:0] kh200=1;	reg signed [w10-1:0] ki200=124;
reg signed [w10-1:0] ka201=-84;	reg signed [w10-1:0] kb201=-34;	reg signed [w10-1:0] kc201=34;	reg signed [w10-1:0] kd201=3;	reg signed [w10-1:0] ke201=-10;	reg signed [w10-1:0] kf201=-110;	reg signed [w10-1:0] kg201=-25;	reg signed [w10-1:0] kh201=90;	reg signed [w10-1:0] ki201=-143;
reg signed [w10-1:0] ka202=-82;	reg signed [w10-1:0] kb202=-50;	reg signed [w10-1:0] kc202=57;	reg signed [w10-1:0] kd202=24;	reg signed [w10-1:0] ke202=-21;	reg signed [w10-1:0] kf202=62;	reg signed [w10-1:0] kg202=89;	reg signed [w10-1:0] kh202=-103;	reg signed [w10-1:0] ki202=90;
reg signed [w10-1:0] ka203=103;	reg signed [w10-1:0] kb203=-22;	reg signed [w10-1:0] kc203=55;	reg signed [w10-1:0] kd203=-107;	reg signed [w10-1:0] ke203=-54;	reg signed [w10-1:0] kf203=120;	reg signed [w10-1:0] kg203=76;	reg signed [w10-1:0] kh203=-114;	reg signed [w10-1:0] ki203=68;
reg signed [w10-1:0] ka204=45;	reg signed [w10-1:0] kb204=-59;	reg signed [w10-1:0] kc204=-40;	reg signed [w10-1:0] kd204=-64;	reg signed [w10-1:0] ke204=-93;	reg signed [w10-1:0] kf204=-61;	reg signed [w10-1:0] kg204=-80;	reg signed [w10-1:0] kh204=-134;	reg signed [w10-1:0] ki204=-70;
reg signed [w10-1:0] ka205=-43;	reg signed [w10-1:0] kb205=-79;	reg signed [w10-1:0] kc205=62;	reg signed [w10-1:0] kd205=-1;	reg signed [w10-1:0] ke205=1;	reg signed [w10-1:0] kf205=-40;	reg signed [w10-1:0] kg205=-107;	reg signed [w10-1:0] kh205=-17;	reg signed [w10-1:0] ki205=55;
reg signed [w10-1:0] ka206=61;	reg signed [w10-1:0] kb206=30;	reg signed [w10-1:0] kc206=-95;	reg signed [w10-1:0] kd206=33;	reg signed [w10-1:0] ke206=-122;	reg signed [w10-1:0] kf206=-88;	reg signed [w10-1:0] kg206=-46;	reg signed [w10-1:0] kh206=35;	reg signed [w10-1:0] ki206=-87;
reg signed [w10-1:0] ka207=-118;	reg signed [w10-1:0] kb207=50;	reg signed [w10-1:0] kc207=-32;	reg signed [w10-1:0] kd207=114;	reg signed [w10-1:0] ke207=25;	reg signed [w10-1:0] kf207=96;	reg signed [w10-1:0] kg207=-6;	reg signed [w10-1:0] kh207=54;	reg signed [w10-1:0] ki207=-15;
reg signed [w10-1:0] ka208=-84;	reg signed [w10-1:0] kb208=-29;	reg signed [w10-1:0] kc208=-101;	reg signed [w10-1:0] kd208=60;	reg signed [w10-1:0] ke208=48;	reg signed [w10-1:0] kf208=31;	reg signed [w10-1:0] kg208=18;	reg signed [w10-1:0] kh208=-32;	reg signed [w10-1:0] ki208=-50;
reg signed [w10-1:0] ka209=-31;	reg signed [w10-1:0] kb209=-106;	reg signed [w10-1:0] kc209=-62;	reg signed [w10-1:0] kd209=9;	reg signed [w10-1:0] ke209=121;	reg signed [w10-1:0] kf209=-125;	reg signed [w10-1:0] kg209=-59;	reg signed [w10-1:0] kh209=-92;	reg signed [w10-1:0] ki209=66;
reg signed [w10-1:0] ka210=-58;	reg signed [w10-1:0] kb210=-22;	reg signed [w10-1:0] kc210=-10;	reg signed [w10-1:0] kd210=78;	reg signed [w10-1:0] ke210=-96;	reg signed [w10-1:0] kf210=-56;	reg signed [w10-1:0] kg210=4;	reg signed [w10-1:0] kh210=-65;	reg signed [w10-1:0] ki210=144;
reg signed [w10-1:0] ka211=-41;	reg signed [w10-1:0] kb211=-42;	reg signed [w10-1:0] kc211=-13;	reg signed [w10-1:0] kd211=111;	reg signed [w10-1:0] ke211=-118;	reg signed [w10-1:0] kf211=-97;	reg signed [w10-1:0] kg211=98;	reg signed [w10-1:0] kh211=-39;	reg signed [w10-1:0] ki211=131;
reg signed [w10-1:0] ka212=-81;	reg signed [w10-1:0] kb212=-13;	reg signed [w10-1:0] kc212=0;	reg signed [w10-1:0] kd212=-82;	reg signed [w10-1:0] ke212=-112;	reg signed [w10-1:0] kf212=91;	reg signed [w10-1:0] kg212=-10;	reg signed [w10-1:0] kh212=-55;	reg signed [w10-1:0] ki212=-42;
reg signed [w10-1:0] ka213=37;	reg signed [w10-1:0] kb213=65;	reg signed [w10-1:0] kc213=5;	reg signed [w10-1:0] kd213=-109;	reg signed [w10-1:0] ke213=-116;	reg signed [w10-1:0] kf213=-45;	reg signed [w10-1:0] kg213=-90;	reg signed [w10-1:0] kh213=-120;	reg signed [w10-1:0] ki213=-88;
reg signed [w10-1:0] ka214=76;	reg signed [w10-1:0] kb214=-35;	reg signed [w10-1:0] kc214=95;	reg signed [w10-1:0] kd214=12;	reg signed [w10-1:0] ke214=-87;	reg signed [w10-1:0] kf214=101;	reg signed [w10-1:0] kg214=-52;	reg signed [w10-1:0] kh214=-56;	reg signed [w10-1:0] ki214=105;
reg signed [w10-1:0] ka215=-68;	reg signed [w10-1:0] kb215=-89;	reg signed [w10-1:0] kc215=80;	reg signed [w10-1:0] kd215=29;	reg signed [w10-1:0] ke215=51;	reg signed [w10-1:0] kf215=83;	reg signed [w10-1:0] kg215=-34;	reg signed [w10-1:0] kh215=98;	reg signed [w10-1:0] ki215=-43;
reg signed [w10-1:0] ka216=6;	reg signed [w10-1:0] kb216=-95;	reg signed [w10-1:0] kc216=-56;	reg signed [w10-1:0] kd216=2;	reg signed [w10-1:0] ke216=-7;	reg signed [w10-1:0] kf216=-47;	reg signed [w10-1:0] kg216=90;	reg signed [w10-1:0] kh216=37;	reg signed [w10-1:0] ki216=-10;
reg signed [w10-1:0] ka217=-25;	reg signed [w10-1:0] kb217=0;	reg signed [w10-1:0] kc217=26;	reg signed [w10-1:0] kd217=-37;	reg signed [w10-1:0] ke217=68;	reg signed [w10-1:0] kf217=-128;	reg signed [w10-1:0] kg217=120;	reg signed [w10-1:0] kh217=-41;	reg signed [w10-1:0] ki217=-14;
reg signed [w10-1:0] ka218=-29;	reg signed [w10-1:0] kb218=-36;	reg signed [w10-1:0] kc218=28;	reg signed [w10-1:0] kd218=47;	reg signed [w10-1:0] ke218=10;	reg signed [w10-1:0] kf218=33;	reg signed [w10-1:0] kg218=68;	reg signed [w10-1:0] kh218=39;	reg signed [w10-1:0] ki218=-106;
reg signed [w10-1:0] ka219=-54;	reg signed [w10-1:0] kb219=16;	reg signed [w10-1:0] kc219=-13;	reg signed [w10-1:0] kd219=-116;	reg signed [w10-1:0] ke219=42;	reg signed [w10-1:0] kf219=70;	reg signed [w10-1:0] kg219=1;	reg signed [w10-1:0] kh219=90;	reg signed [w10-1:0] ki219=-5;
reg signed [w10-1:0] ka220=-104;	reg signed [w10-1:0] kb220=-56;	reg signed [w10-1:0] kc220=75;	reg signed [w10-1:0] kd220=43;	reg signed [w10-1:0] ke220=-100;	reg signed [w10-1:0] kf220=-74;	reg signed [w10-1:0] kg220=-12;	reg signed [w10-1:0] kh220=-36;	reg signed [w10-1:0] ki220=-63;
reg signed [w10-1:0] ka221=-34;	reg signed [w10-1:0] kb221=-49;	reg signed [w10-1:0] kc221=-16;	reg signed [w10-1:0] kd221=-14;	reg signed [w10-1:0] ke221=-78;	reg signed [w10-1:0] kf221=96;	reg signed [w10-1:0] kg221=53;	reg signed [w10-1:0] kh221=-45;	reg signed [w10-1:0] ki221=-86;
reg signed [w10-1:0] ka222=60;	reg signed [w10-1:0] kb222=-175;	reg signed [w10-1:0] kc222=1;	reg signed [w10-1:0] kd222=73;	reg signed [w10-1:0] ke222=-21;	reg signed [w10-1:0] kf222=89;	reg signed [w10-1:0] kg222=-51;	reg signed [w10-1:0] kh222=44;	reg signed [w10-1:0] ki222=85;
reg signed [w10-1:0] ka223=148;	reg signed [w10-1:0] kb223=-92;	reg signed [w10-1:0] kc223=81;	reg signed [w10-1:0] kd223=-109;	reg signed [w10-1:0] ke223=-17;	reg signed [w10-1:0] kf223=-36;	reg signed [w10-1:0] kg223=65;	reg signed [w10-1:0] kh223=9;	reg signed [w10-1:0] ki223=30;
reg signed [w10-1:0] ka224=112;	reg signed [w10-1:0] kb224=-17;	reg signed [w10-1:0] kc224=61;	reg signed [w10-1:0] kd224=55;	reg signed [w10-1:0] ke224=-58;	reg signed [w10-1:0] kf224=56;	reg signed [w10-1:0] kg224=125;	reg signed [w10-1:0] kh224=103;	reg signed [w10-1:0] ki224=-153;
reg signed [w10-1:0] ka225=-63;	reg signed [w10-1:0] kb225=-35;	reg signed [w10-1:0] kc225=69;	reg signed [w10-1:0] kd225=85;	reg signed [w10-1:0] ke225=61;	reg signed [w10-1:0] kf225=91;	reg signed [w10-1:0] kg225=65;	reg signed [w10-1:0] kh225=11;	reg signed [w10-1:0] ki225=46;
reg signed [w10-1:0] ka226=-48;	reg signed [w10-1:0] kb226=-12;	reg signed [w10-1:0] kc226=-15;	reg signed [w10-1:0] kd226=-95;	reg signed [w10-1:0] ke226=-95;	reg signed [w10-1:0] kf226=-7;	reg signed [w10-1:0] kg226=-137;	reg signed [w10-1:0] kh226=-91;	reg signed [w10-1:0] ki226=-76;
reg signed [w10-1:0] ka227=44;	reg signed [w10-1:0] kb227=55;	reg signed [w10-1:0] kc227=38;	reg signed [w10-1:0] kd227=-95;	reg signed [w10-1:0] ke227=-45;	reg signed [w10-1:0] kf227=90;	reg signed [w10-1:0] kg227=-84;	reg signed [w10-1:0] kh227=-37;	reg signed [w10-1:0] ki227=120;
reg signed [w10-1:0] ka228=34;	reg signed [w10-1:0] kb228=52;	reg signed [w10-1:0] kc228=68;	reg signed [w10-1:0] kd228=-21;	reg signed [w10-1:0] ke228=4;	reg signed [w10-1:0] kf228=-67;	reg signed [w10-1:0] kg228=-31;	reg signed [w10-1:0] kh228=-103;	reg signed [w10-1:0] ki228=-99;
reg signed [w10-1:0] ka229=-20;	reg signed [w10-1:0] kb229=76;	reg signed [w10-1:0] kc229=-97;	reg signed [w10-1:0] kd229=-85;	reg signed [w10-1:0] ke229=35;	reg signed [w10-1:0] kf229=76;	reg signed [w10-1:0] kg229=34;	reg signed [w10-1:0] kh229=-126;	reg signed [w10-1:0] ki229=-39;
reg signed [w10-1:0] ka230=121;	reg signed [w10-1:0] kb230=-130;	reg signed [w10-1:0] kc230=77;	reg signed [w10-1:0] kd230=-132;	reg signed [w10-1:0] ke230=-27;	reg signed [w10-1:0] kf230=111;	reg signed [w10-1:0] kg230=7;	reg signed [w10-1:0] kh230=-18;	reg signed [w10-1:0] ki230=11;
reg signed [w10-1:0] ka231=96;	reg signed [w10-1:0] kb231=46;	reg signed [w10-1:0] kc231=-76;	reg signed [w10-1:0] kd231=-71;	reg signed [w10-1:0] ke231=23;	reg signed [w10-1:0] kf231=68;	reg signed [w10-1:0] kg231=-85;	reg signed [w10-1:0] kh231=21;	reg signed [w10-1:0] ki231=89;
reg signed [w10-1:0] ka232=-79;	reg signed [w10-1:0] kb232=-5;	reg signed [w10-1:0] kc232=31;	reg signed [w10-1:0] kd232=38;	reg signed [w10-1:0] ke232=108;	reg signed [w10-1:0] kf232=-67;	reg signed [w10-1:0] kg232=154;	reg signed [w10-1:0] kh232=19;	reg signed [w10-1:0] ki232=-16;
reg signed [w10-1:0] ka233=173;	reg signed [w10-1:0] kb233=-39;	reg signed [w10-1:0] kc233=-1;	reg signed [w10-1:0] kd233=108;	reg signed [w10-1:0] ke233=-128;	reg signed [w10-1:0] kf233=45;	reg signed [w10-1:0] kg233=-21;	reg signed [w10-1:0] kh233=-53;	reg signed [w10-1:0] ki233=-7;
reg signed [w10-1:0] ka234=102;	reg signed [w10-1:0] kb234=125;	reg signed [w10-1:0] kc234=50;	reg signed [w10-1:0] kd234=51;	reg signed [w10-1:0] ke234=-35;	reg signed [w10-1:0] kf234=66;	reg signed [w10-1:0] kg234=-101;	reg signed [w10-1:0] kh234=8;	reg signed [w10-1:0] ki234=-44;
reg signed [w10-1:0] ka235=25;	reg signed [w10-1:0] kb235=9;	reg signed [w10-1:0] kc235=65;	reg signed [w10-1:0] kd235=-72;	reg signed [w10-1:0] ke235=-67;	reg signed [w10-1:0] kf235=1;	reg signed [w10-1:0] kg235=-20;	reg signed [w10-1:0] kh235=29;	reg signed [w10-1:0] ki235=-97;
reg signed [w10-1:0] ka236=-60;	reg signed [w10-1:0] kb236=-117;	reg signed [w10-1:0] kc236=-40;	reg signed [w10-1:0] kd236=-91;	reg signed [w10-1:0] ke236=49;	reg signed [w10-1:0] kf236=65;	reg signed [w10-1:0] kg236=-97;	reg signed [w10-1:0] kh236=8;	reg signed [w10-1:0] ki236=34;
reg signed [w10-1:0] ka237=94;	reg signed [w10-1:0] kb237=60;	reg signed [w10-1:0] kc237=75;	reg signed [w10-1:0] kd237=4;	reg signed [w10-1:0] ke237=38;	reg signed [w10-1:0] kf237=-99;	reg signed [w10-1:0] kg237=-17;	reg signed [w10-1:0] kh237=48;	reg signed [w10-1:0] ki237=-7;
reg signed [w10-1:0] ka238=-37;	reg signed [w10-1:0] kb238=24;	reg signed [w10-1:0] kc238=47;	reg signed [w10-1:0] kd238=1;	reg signed [w10-1:0] ke238=-91;	reg signed [w10-1:0] kf238=48;	reg signed [w10-1:0] kg238=-80;	reg signed [w10-1:0] kh238=-2;	reg signed [w10-1:0] ki238=-19;
reg signed [w10-1:0] ka239=-164;	reg signed [w10-1:0] kb239=122;	reg signed [w10-1:0] kc239=144;	reg signed [w10-1:0] kd239=-113;	reg signed [w10-1:0] ke239=72;	reg signed [w10-1:0] kf239=94;	reg signed [w10-1:0] kg239=-98;	reg signed [w10-1:0] kh239=-43;	reg signed [w10-1:0] ki239=4;
reg signed [w10-1:0] ka240=-118;	reg signed [w10-1:0] kb240=13;	reg signed [w10-1:0] kc240=85;	reg signed [w10-1:0] kd240=-63;	reg signed [w10-1:0] ke240=108;	reg signed [w10-1:0] kf240=-134;	reg signed [w10-1:0] kg240=78;	reg signed [w10-1:0] kh240=-82;	reg signed [w10-1:0] ki240=22;
reg signed [w10-1:0] ka241=-117;	reg signed [w10-1:0] kb241=-61;	reg signed [w10-1:0] kc241=-40;	reg signed [w10-1:0] kd241=76;	reg signed [w10-1:0] ke241=-13;	reg signed [w10-1:0] kf241=-120;	reg signed [w10-1:0] kg241=6;	reg signed [w10-1:0] kh241=70;	reg signed [w10-1:0] ki241=6;
reg signed [w10-1:0] ka242=-34;	reg signed [w10-1:0] kb242=-27;	reg signed [w10-1:0] kc242=56;	reg signed [w10-1:0] kd242=-105;	reg signed [w10-1:0] ke242=-63;	reg signed [w10-1:0] kf242=-87;	reg signed [w10-1:0] kg242=35;	reg signed [w10-1:0] kh242=90;	reg signed [w10-1:0] ki242=2;
reg signed [w10-1:0] ka243=116;	reg signed [w10-1:0] kb243=21;	reg signed [w10-1:0] kc243=115;	reg signed [w10-1:0] kd243=-25;	reg signed [w10-1:0] ke243=9;	reg signed [w10-1:0] kf243=124;	reg signed [w10-1:0] kg243=61;	reg signed [w10-1:0] kh243=-102;	reg signed [w10-1:0] ki243=9;
reg signed [w10-1:0] ka244=-14;	reg signed [w10-1:0] kb244=-85;	reg signed [w10-1:0] kc244=-79;	reg signed [w10-1:0] kd244=93;	reg signed [w10-1:0] ke244=46;	reg signed [w10-1:0] kf244=-173;	reg signed [w10-1:0] kg244=-17;	reg signed [w10-1:0] kh244=9;	reg signed [w10-1:0] ki244=-82;
reg signed [w10-1:0] ka245=-107;	reg signed [w10-1:0] kb245=-115;	reg signed [w10-1:0] kc245=-11;	reg signed [w10-1:0] kd245=80;	reg signed [w10-1:0] ke245=-27;	reg signed [w10-1:0] kf245=12;	reg signed [w10-1:0] kg245=108;	reg signed [w10-1:0] kh245=28;	reg signed [w10-1:0] ki245=-36;
reg signed [w10-1:0] ka246=-51;	reg signed [w10-1:0] kb246=-12;	reg signed [w10-1:0] kc246=-122;	reg signed [w10-1:0] kd246=-49;	reg signed [w10-1:0] ke246=-25;	reg signed [w10-1:0] kf246=-56;	reg signed [w10-1:0] kg246=71;	reg signed [w10-1:0] kh246=46;	reg signed [w10-1:0] ki246=34;
reg signed [w10-1:0] ka247=110;	reg signed [w10-1:0] kb247=-29;	reg signed [w10-1:0] kc247=107;	reg signed [w10-1:0] kd247=-4;	reg signed [w10-1:0] ke247=-14;	reg signed [w10-1:0] kf247=-39;	reg signed [w10-1:0] kg247=19;	reg signed [w10-1:0] kh247=-64;	reg signed [w10-1:0] ki247=100;
reg signed [w10-1:0] ka248=-94;	reg signed [w10-1:0] kb248=72;	reg signed [w10-1:0] kc248=-39;	reg signed [w10-1:0] kd248=41;	reg signed [w10-1:0] ke248=32;	reg signed [w10-1:0] kf248=-76;	reg signed [w10-1:0] kg248=-34;	reg signed [w10-1:0] kh248=-128;	reg signed [w10-1:0] ki248=53;
reg signed [w10-1:0] ka249=-16;	reg signed [w10-1:0] kb249=-100;	reg signed [w10-1:0] kc249=43;	reg signed [w10-1:0] kd249=-51;	reg signed [w10-1:0] ke249=-22;	reg signed [w10-1:0] kf249=15;	reg signed [w10-1:0] kg249=-52;	reg signed [w10-1:0] kh249=-20;	reg signed [w10-1:0] ki249=84;
reg signed [w10-1:0] ka250=9;	reg signed [w10-1:0] kb250=145;	reg signed [w10-1:0] kc250=66;	reg signed [w10-1:0] kd250=68;	reg signed [w10-1:0] ke250=64;	reg signed [w10-1:0] kf250=114;	reg signed [w10-1:0] kg250=-30;	reg signed [w10-1:0] kh250=-105;	reg signed [w10-1:0] ki250=-52;
reg signed [w10-1:0] ka251=-84;	reg signed [w10-1:0] kb251=18;	reg signed [w10-1:0] kc251=-110;	reg signed [w10-1:0] kd251=42;	reg signed [w10-1:0] ke251=57;	reg signed [w10-1:0] kf251=-28;	reg signed [w10-1:0] kg251=-97;	reg signed [w10-1:0] kh251=-15;	reg signed [w10-1:0] ki251=68;
reg signed [w10-1:0] ka252=-43;	reg signed [w10-1:0] kb252=-54;	reg signed [w10-1:0] kc252=103;	reg signed [w10-1:0] kd252=74;	reg signed [w10-1:0] ke252=-116;	reg signed [w10-1:0] kf252=75;	reg signed [w10-1:0] kg252=-31;	reg signed [w10-1:0] kh252=100;	reg signed [w10-1:0] ki252=-93;
reg signed [w10-1:0] ka253=91;	reg signed [w10-1:0] kb253=110;	reg signed [w10-1:0] kc253=-91;	reg signed [w10-1:0] kd253=18;	reg signed [w10-1:0] ke253=-63;	reg signed [w10-1:0] kf253=-87;	reg signed [w10-1:0] kg253=44;	reg signed [w10-1:0] kh253=34;	reg signed [w10-1:0] ki253=60;
reg signed [w10-1:0] ka254=37;	reg signed [w10-1:0] kb254=70;	reg signed [w10-1:0] kc254=-75;	reg signed [w10-1:0] kd254=57;	reg signed [w10-1:0] ke254=-48;	reg signed [w10-1:0] kf254=51;	reg signed [w10-1:0] kg254=-63;	reg signed [w10-1:0] kh254=-9;	reg signed [w10-1:0] ki254=106;
reg signed [w10-1:0] ka255=59;	reg signed [w10-1:0] kb255=-131;	reg signed [w10-1:0] kc255=56;	reg signed [w10-1:0] kd255=-66;	reg signed [w10-1:0] ke255=-25;	reg signed [w10-1:0] kf255=-67;	reg signed [w10-1:0] kg255=-3;	reg signed [w10-1:0] kh255=144;	reg signed [w10-1:0] ki255=-13;
reg signed [w10-1:0] ka256=31;	reg signed [w10-1:0] kb256=-40;	reg signed [w10-1:0] kc256=12;	reg signed [w10-1:0] kd256=5;	reg signed [w10-1:0] ke256=-37;	reg signed [w10-1:0] kf256=37;	reg signed [w10-1:0] kg256=-86;	reg signed [w10-1:0] kh256=-102;	reg signed [w10-1:0] ki256=78;
reg signed [w10-1:0] ka257=8;	reg signed [w10-1:0] kb257=-44;	reg signed [w10-1:0] kc257=-10;	reg signed [w10-1:0] kd257=76;	reg signed [w10-1:0] ke257=49;	reg signed [w10-1:0] kf257=-27;	reg signed [w10-1:0] kg257=108;	reg signed [w10-1:0] kh257=121;	reg signed [w10-1:0] ki257=-38;
reg signed [w10-1:0] ka258=-49;	reg signed [w10-1:0] kb258=-79;	reg signed [w10-1:0] kc258=-85;	reg signed [w10-1:0] kd258=98;	reg signed [w10-1:0] ke258=-33;	reg signed [w10-1:0] kf258=20;	reg signed [w10-1:0] kg258=16;	reg signed [w10-1:0] kh258=78;	reg signed [w10-1:0] ki258=-11;
reg signed [w10-1:0] ka259=35;	reg signed [w10-1:0] kb259=-22;	reg signed [w10-1:0] kc259=6;	reg signed [w10-1:0] kd259=-115;	reg signed [w10-1:0] ke259=6;	reg signed [w10-1:0] kf259=-95;	reg signed [w10-1:0] kg259=70;	reg signed [w10-1:0] kh259=-122;	reg signed [w10-1:0] ki259=-83;
reg signed [w10-1:0] ka260=-102;	reg signed [w10-1:0] kb260=15;	reg signed [w10-1:0] kc260=-102;	reg signed [w10-1:0] kd260=14;	reg signed [w10-1:0] ke260=107;	reg signed [w10-1:0] kf260=-82;	reg signed [w10-1:0] kg260=59;	reg signed [w10-1:0] kh260=13;	reg signed [w10-1:0] ki260=60;
reg signed [w10-1:0] ka261=68;	reg signed [w10-1:0] kb261=118;	reg signed [w10-1:0] kc261=-1;	reg signed [w10-1:0] kd261=94;	reg signed [w10-1:0] ke261=-13;	reg signed [w10-1:0] kf261=20;	reg signed [w10-1:0] kg261=-57;	reg signed [w10-1:0] kh261=54;	reg signed [w10-1:0] ki261=-63;
reg signed [w10-1:0] ka262=24;	reg signed [w10-1:0] kb262=-30;	reg signed [w10-1:0] kc262=99;	reg signed [w10-1:0] kd262=-73;	reg signed [w10-1:0] ke262=-35;	reg signed [w10-1:0] kf262=-69;	reg signed [w10-1:0] kg262=-128;	reg signed [w10-1:0] kh262=-159;	reg signed [w10-1:0] ki262=102;
reg signed [w10-1:0] ka263=-141;	reg signed [w10-1:0] kb263=-44;	reg signed [w10-1:0] kc263=-99;	reg signed [w10-1:0] kd263=-60;	reg signed [w10-1:0] ke263=55;	reg signed [w10-1:0] kf263=-108;	reg signed [w10-1:0] kg263=-76;	reg signed [w10-1:0] kh263=-41;	reg signed [w10-1:0] ki263=-26;
reg signed [w10-1:0] ka264=56;	reg signed [w10-1:0] kb264=49;	reg signed [w10-1:0] kc264=10;	reg signed [w10-1:0] kd264=-9;	reg signed [w10-1:0] ke264=66;	reg signed [w10-1:0] kf264=46;	reg signed [w10-1:0] kg264=127;	reg signed [w10-1:0] kh264=-41;	reg signed [w10-1:0] ki264=33;
reg signed [w10-1:0] ka265=39;	reg signed [w10-1:0] kb265=-91;	reg signed [w10-1:0] kc265=-60;	reg signed [w10-1:0] kd265=-52;	reg signed [w10-1:0] ke265=-10;	reg signed [w10-1:0] kf265=-13;	reg signed [w10-1:0] kg265=152;	reg signed [w10-1:0] kh265=136;	reg signed [w10-1:0] ki265=-97;
reg signed [w10-1:0] ka266=62;	reg signed [w10-1:0] kb266=-24;	reg signed [w10-1:0] kc266=-86;	reg signed [w10-1:0] kd266=54;	reg signed [w10-1:0] ke266=-48;	reg signed [w10-1:0] kf266=-6;	reg signed [w10-1:0] kg266=-66;	reg signed [w10-1:0] kh266=-113;	reg signed [w10-1:0] ki266=5;
reg signed [w10-1:0] ka267=97;	reg signed [w10-1:0] kb267=113;	reg signed [w10-1:0] kc267=31;	reg signed [w10-1:0] kd267=-23;	reg signed [w10-1:0] ke267=-37;	reg signed [w10-1:0] kf267=97;	reg signed [w10-1:0] kg267=-7;	reg signed [w10-1:0] kh267=-73;	reg signed [w10-1:0] ki267=-7;
reg signed [w10-1:0] ka268=-24;	reg signed [w10-1:0] kb268=30;	reg signed [w10-1:0] kc268=60;	reg signed [w10-1:0] kd268=-108;	reg signed [w10-1:0] ke268=41;	reg signed [w10-1:0] kf268=53;	reg signed [w10-1:0] kg268=-55;	reg signed [w10-1:0] kh268=92;	reg signed [w10-1:0] ki268=-99;
reg signed [w10-1:0] ka269=46;	reg signed [w10-1:0] kb269=37;	reg signed [w10-1:0] kc269=54;	reg signed [w10-1:0] kd269=-115;	reg signed [w10-1:0] ke269=-79;	reg signed [w10-1:0] kf269=30;	reg signed [w10-1:0] kg269=50;	reg signed [w10-1:0] kh269=110;	reg signed [w10-1:0] ki269=5;
reg signed [w10-1:0] ka270=34;	reg signed [w10-1:0] kb270=138;	reg signed [w10-1:0] kc270=98;	reg signed [w10-1:0] kd270=-8;	reg signed [w10-1:0] ke270=30;	reg signed [w10-1:0] kf270=-13;	reg signed [w10-1:0] kg270=-51;	reg signed [w10-1:0] kh270=-110;	reg signed [w10-1:0] ki270=-55;
reg signed [w10-1:0] ka271=-74;	reg signed [w10-1:0] kb271=-130;	reg signed [w10-1:0] kc271=28;	reg signed [w10-1:0] kd271=67;	reg signed [w10-1:0] ke271=-76;	reg signed [w10-1:0] kf271=-37;	reg signed [w10-1:0] kg271=58;	reg signed [w10-1:0] kh271=93;	reg signed [w10-1:0] ki271=-60;
reg signed [w10-1:0] ka272=-87;	reg signed [w10-1:0] kb272=-12;	reg signed [w10-1:0] kc272=-76;	reg signed [w10-1:0] kd272=-16;	reg signed [w10-1:0] ke272=-29;	reg signed [w10-1:0] kf272=52;	reg signed [w10-1:0] kg272=-103;	reg signed [w10-1:0] kh272=-42;	reg signed [w10-1:0] ki272=-70;
reg signed [w10-1:0] ka273=19;	reg signed [w10-1:0] kb273=60;	reg signed [w10-1:0] kc273=52;	reg signed [w10-1:0] kd273=-60;	reg signed [w10-1:0] ke273=-97;	reg signed [w10-1:0] kf273=136;	reg signed [w10-1:0] kg273=-22;	reg signed [w10-1:0] kh273=90;	reg signed [w10-1:0] ki273=-70;
reg signed [w10-1:0] ka274=1;	reg signed [w10-1:0] kb274=14;	reg signed [w10-1:0] kc274=34;	reg signed [w10-1:0] kd274=65;	reg signed [w10-1:0] ke274=125;	reg signed [w10-1:0] kf274=48;	reg signed [w10-1:0] kg274=67;	reg signed [w10-1:0] kh274=-120;	reg signed [w10-1:0] ki274=79;
reg signed [w10-1:0] ka275=-41;	reg signed [w10-1:0] kb275=-87;	reg signed [w10-1:0] kc275=13;	reg signed [w10-1:0] kd275=27;	reg signed [w10-1:0] ke275=91;	reg signed [w10-1:0] kf275=-63;	reg signed [w10-1:0] kg275=2;	reg signed [w10-1:0] kh275=-107;	reg signed [w10-1:0] ki275=86;
reg signed [w10-1:0] ka276=-22;	reg signed [w10-1:0] kb276=-133;	reg signed [w10-1:0] kc276=49;	reg signed [w10-1:0] kd276=-81;	reg signed [w10-1:0] ke276=-52;	reg signed [w10-1:0] kf276=-52;	reg signed [w10-1:0] kg276=137;	reg signed [w10-1:0] kh276=-15;	reg signed [w10-1:0] ki276=-61;
reg signed [w10-1:0] ka277=38;	reg signed [w10-1:0] kb277=90;	reg signed [w10-1:0] kc277=116;	reg signed [w10-1:0] kd277=-26;	reg signed [w10-1:0] ke277=26;	reg signed [w10-1:0] kf277=-97;	reg signed [w10-1:0] kg277=151;	reg signed [w10-1:0] kh277=58;	reg signed [w10-1:0] ki277=-61;
reg signed [w10-1:0] ka278=-100;	reg signed [w10-1:0] kb278=161;	reg signed [w10-1:0] kc278=25;	reg signed [w10-1:0] kd278=-39;	reg signed [w10-1:0] ke278=6;	reg signed [w10-1:0] kf278=48;	reg signed [w10-1:0] kg278=-108;	reg signed [w10-1:0] kh278=42;	reg signed [w10-1:0] ki278=87;
reg signed [w10-1:0] ka279=-43;	reg signed [w10-1:0] kb279=10;	reg signed [w10-1:0] kc279=-2;	reg signed [w10-1:0] kd279=-44;	reg signed [w10-1:0] ke279=13;	reg signed [w10-1:0] kf279=-25;	reg signed [w10-1:0] kg279=-105;	reg signed [w10-1:0] kh279=26;	reg signed [w10-1:0] ki279=-117;
reg signed [w10-1:0] ka280=70;	reg signed [w10-1:0] kb280=48;	reg signed [w10-1:0] kc280=-16;	reg signed [w10-1:0] kd280=78;	reg signed [w10-1:0] ke280=74;	reg signed [w10-1:0] kf280=22;	reg signed [w10-1:0] kg280=-78;	reg signed [w10-1:0] kh280=-93;	reg signed [w10-1:0] ki280=71;
reg signed [w10-1:0] ka281=130;	reg signed [w10-1:0] kb281=-37;	reg signed [w10-1:0] kc281=-2;	reg signed [w10-1:0] kd281=-12;	reg signed [w10-1:0] ke281=8;	reg signed [w10-1:0] kf281=85;	reg signed [w10-1:0] kg281=5;	reg signed [w10-1:0] kh281=-133;	reg signed [w10-1:0] ki281=63;
reg signed [w10-1:0] ka282=-111;	reg signed [w10-1:0] kb282=108;	reg signed [w10-1:0] kc282=-78;	reg signed [w10-1:0] kd282=114;	reg signed [w10-1:0] ke282=31;	reg signed [w10-1:0] kf282=33;	reg signed [w10-1:0] kg282=-93;	reg signed [w10-1:0] kh282=-96;	reg signed [w10-1:0] ki282=47;
reg signed [w10-1:0] ka283=-122;	reg signed [w10-1:0] kb283=19;	reg signed [w10-1:0] kc283=72;	reg signed [w10-1:0] kd283=-65;	reg signed [w10-1:0] ke283=83;	reg signed [w10-1:0] kf283=11;	reg signed [w10-1:0] kg283=-75;	reg signed [w10-1:0] kh283=15;	reg signed [w10-1:0] ki283=121;
reg signed [w10-1:0] ka284=-72;	reg signed [w10-1:0] kb284=-127;	reg signed [w10-1:0] kc284=60;	reg signed [w10-1:0] kd284=65;	reg signed [w10-1:0] ke284=-105;	reg signed [w10-1:0] kf284=-147;	reg signed [w10-1:0] kg284=13;	reg signed [w10-1:0] kh284=30;	reg signed [w10-1:0] ki284=-6;
reg signed [w10-1:0] ka285=76;	reg signed [w10-1:0] kb285=14;	reg signed [w10-1:0] kc285=-29;	reg signed [w10-1:0] kd285=117;	reg signed [w10-1:0] ke285=-27;	reg signed [w10-1:0] kf285=56;	reg signed [w10-1:0] kg285=126;	reg signed [w10-1:0] kh285=-19;	reg signed [w10-1:0] ki285=57;
reg signed [w10-1:0] ka286=82;	reg signed [w10-1:0] kb286=90;	reg signed [w10-1:0] kc286=91;	reg signed [w10-1:0] kd286=-96;	reg signed [w10-1:0] ke286=-104;	reg signed [w10-1:0] kf286=-77;	reg signed [w10-1:0] kg286=-41;	reg signed [w10-1:0] kh286=-48;	reg signed [w10-1:0] ki286=-56;
reg signed [w10-1:0] ka287=6;	reg signed [w10-1:0] kb287=-5;	reg signed [w10-1:0] kc287=-134;	reg signed [w10-1:0] kd287=-32;	reg signed [w10-1:0] ke287=-88;	reg signed [w10-1:0] kf287=3;	reg signed [w10-1:0] kg287=-78;	reg signed [w10-1:0] kh287=11;	reg signed [w10-1:0] ki287=14;
reg signed [w10-1:0] ka288=50;	reg signed [w10-1:0] kb288=1;	reg signed [w10-1:0] kc288=-14;	reg signed [w10-1:0] kd288=-26;	reg signed [w10-1:0] ke288=20;	reg signed [w10-1:0] kf288=-36;	reg signed [w10-1:0] kg288=-30;	reg signed [w10-1:0] kh288=-95;	reg signed [w10-1:0] ki288=-83;
reg signed [w10-1:0] ka289=-43;	reg signed [w10-1:0] kb289=29;	reg signed [w10-1:0] kc289=54;	reg signed [w10-1:0] kd289=-54;	reg signed [w10-1:0] ke289=16;	reg signed [w10-1:0] kf289=42;	reg signed [w10-1:0] kg289=46;	reg signed [w10-1:0] kh289=94;	reg signed [w10-1:0] ki289=-34;
reg signed [w10-1:0] ka290=-117;	reg signed [w10-1:0] kb290=47;	reg signed [w10-1:0] kc290=51;	reg signed [w10-1:0] kd290=101;	reg signed [w10-1:0] ke290=-125;	reg signed [w10-1:0] kf290=70;	reg signed [w10-1:0] kg290=42;	reg signed [w10-1:0] kh290=56;	reg signed [w10-1:0] ki290=18;
reg signed [w10-1:0] ka291=-56;	reg signed [w10-1:0] kb291=-48;	reg signed [w10-1:0] kc291=-121;	reg signed [w10-1:0] kd291=-100;	reg signed [w10-1:0] ke291=86;	reg signed [w10-1:0] kf291=-52;	reg signed [w10-1:0] kg291=-22;	reg signed [w10-1:0] kh291=127;	reg signed [w10-1:0] ki291=153;
reg signed [w10-1:0] ka292=15;	reg signed [w10-1:0] kb292=-3;	reg signed [w10-1:0] kc292=18;	reg signed [w10-1:0] kd292=16;	reg signed [w10-1:0] ke292=-82;	reg signed [w10-1:0] kf292=-4;	reg signed [w10-1:0] kg292=-59;	reg signed [w10-1:0] kh292=-20;	reg signed [w10-1:0] ki292=-74;
reg signed [w10-1:0] ka293=54;	reg signed [w10-1:0] kb293=-33;	reg signed [w10-1:0] kc293=-74;	reg signed [w10-1:0] kd293=-69;	reg signed [w10-1:0] ke293=-106;	reg signed [w10-1:0] kf293=-53;	reg signed [w10-1:0] kg293=-15;	reg signed [w10-1:0] kh293=-59;	reg signed [w10-1:0] ki293=-14;
reg signed [w10-1:0] ka294=85;	reg signed [w10-1:0] kb294=142;	reg signed [w10-1:0] kc294=42;	reg signed [w10-1:0] kd294=81;	reg signed [w10-1:0] ke294=55;	reg signed [w10-1:0] kf294=-89;	reg signed [w10-1:0] kg294=-74;	reg signed [w10-1:0] kh294=64;	reg signed [w10-1:0] ki294=110;
reg signed [w10-1:0] ka295=4;	reg signed [w10-1:0] kb295=-38;	reg signed [w10-1:0] kc295=-128;	reg signed [w10-1:0] kd295=-88;	reg signed [w10-1:0] ke295=139;	reg signed [w10-1:0] kf295=99;	reg signed [w10-1:0] kg295=90;	reg signed [w10-1:0] kh295=-77;	reg signed [w10-1:0] ki295=92;
reg signed [w10-1:0] ka296=-5;	reg signed [w10-1:0] kb296=35;	reg signed [w10-1:0] kc296=26;	reg signed [w10-1:0] kd296=-75;	reg signed [w10-1:0] ke296=132;	reg signed [w10-1:0] kf296=88;	reg signed [w10-1:0] kg296=27;	reg signed [w10-1:0] kh296=131;	reg signed [w10-1:0] ki296=-84;
reg signed [w10-1:0] ka297=-80;	reg signed [w10-1:0] kb297=67;	reg signed [w10-1:0] kc297=9;	reg signed [w10-1:0] kd297=-171;	reg signed [w10-1:0] ke297=-43;	reg signed [w10-1:0] kf297=-87;	reg signed [w10-1:0] kg297=-138;	reg signed [w10-1:0] kh297=41;	reg signed [w10-1:0] ki297=-64;
reg signed [w10-1:0] ka298=-56;	reg signed [w10-1:0] kb298=101;	reg signed [w10-1:0] kc298=-88;	reg signed [w10-1:0] kd298=4;	reg signed [w10-1:0] ke298=-97;	reg signed [w10-1:0] kf298=44;	reg signed [w10-1:0] kg298=-76;	reg signed [w10-1:0] kh298=90;	reg signed [w10-1:0] ki298=-82;
reg signed [w10-1:0] ka299=35;	reg signed [w10-1:0] kb299=-37;	reg signed [w10-1:0] kc299=-40;	reg signed [w10-1:0] kd299=-43;	reg signed [w10-1:0] ke299=5;	reg signed [w10-1:0] kf299=-28;	reg signed [w10-1:0] kg299=172;	reg signed [w10-1:0] kh299=-26;	reg signed [w10-1:0] ki299=25;
reg signed [w10-1:0] ka300=32;	reg signed [w10-1:0] kb300=33;	reg signed [w10-1:0] kc300=99;	reg signed [w10-1:0] kd300=-98;	reg signed [w10-1:0] ke300=19;	reg signed [w10-1:0] kf300=-25;	reg signed [w10-1:0] kg300=-37;	reg signed [w10-1:0] kh300=-124;	reg signed [w10-1:0] ki300=101;
reg signed [w10-1:0] ka301=-39;	reg signed [w10-1:0] kb301=50;	reg signed [w10-1:0] kc301=66;	reg signed [w10-1:0] kd301=106;	reg signed [w10-1:0] ke301=-102;	reg signed [w10-1:0] kf301=-5;	reg signed [w10-1:0] kg301=33;	reg signed [w10-1:0] kh301=59;	reg signed [w10-1:0] ki301=16;
reg signed [w10-1:0] ka302=36;	reg signed [w10-1:0] kb302=4;	reg signed [w10-1:0] kc302=-76;	reg signed [w10-1:0] kd302=-34;	reg signed [w10-1:0] ke302=21;	reg signed [w10-1:0] kf302=-38;	reg signed [w10-1:0] kg302=-31;	reg signed [w10-1:0] kh302=5;	reg signed [w10-1:0] ki302=135;
reg signed [w10-1:0] ka303=-6;	reg signed [w10-1:0] kb303=-74;	reg signed [w10-1:0] kc303=24;	reg signed [w10-1:0] kd303=29;	reg signed [w10-1:0] ke303=119;	reg signed [w10-1:0] kf303=83;	reg signed [w10-1:0] kg303=91;	reg signed [w10-1:0] kh303=29;	reg signed [w10-1:0] ki303=-42;
reg signed [w10-1:0] ka304=120;	reg signed [w10-1:0] kb304=-47;	reg signed [w10-1:0] kc304=-20;	reg signed [w10-1:0] kd304=-35;	reg signed [w10-1:0] ke304=139;	reg signed [w10-1:0] kf304=-40;	reg signed [w10-1:0] kg304=-17;	reg signed [w10-1:0] kh304=21;	reg signed [w10-1:0] ki304=-99;
reg signed [w10-1:0] ka305=32;	reg signed [w10-1:0] kb305=171;	reg signed [w10-1:0] kc305=56;	reg signed [w10-1:0] kd305=-37;	reg signed [w10-1:0] ke305=122;	reg signed [w10-1:0] kf305=22;	reg signed [w10-1:0] kg305=16;	reg signed [w10-1:0] kh305=163;	reg signed [w10-1:0] ki305=-12;
reg signed [w10-1:0] ka306=27;	reg signed [w10-1:0] kb306=54;	reg signed [w10-1:0] kc306=37;	reg signed [w10-1:0] kd306=-108;	reg signed [w10-1:0] ke306=31;	reg signed [w10-1:0] kf306=-27;	reg signed [w10-1:0] kg306=-66;	reg signed [w10-1:0] kh306=-17;	reg signed [w10-1:0] ki306=-57;
reg signed [w10-1:0] ka307=-40;	reg signed [w10-1:0] kb307=34;	reg signed [w10-1:0] kc307=40;	reg signed [w10-1:0] kd307=-124;	reg signed [w10-1:0] ke307=4;	reg signed [w10-1:0] kf307=-12;	reg signed [w10-1:0] kg307=74;	reg signed [w10-1:0] kh307=66;	reg signed [w10-1:0] ki307=1;
reg signed [w10-1:0] ka308=197;	reg signed [w10-1:0] kb308=52;	reg signed [w10-1:0] kc308=21;	reg signed [w10-1:0] kd308=32;	reg signed [w10-1:0] ke308=-102;	reg signed [w10-1:0] kf308=-63;	reg signed [w10-1:0] kg308=67;	reg signed [w10-1:0] kh308=-5;	reg signed [w10-1:0] ki308=13;
reg signed [w10-1:0] ka309=-63;	reg signed [w10-1:0] kb309=-53;	reg signed [w10-1:0] kc309=103;	reg signed [w10-1:0] kd309=-48;	reg signed [w10-1:0] ke309=-7;	reg signed [w10-1:0] kf309=102;	reg signed [w10-1:0] kg309=-95;	reg signed [w10-1:0] kh309=22;	reg signed [w10-1:0] ki309=-58;
reg signed [w10-1:0] ka310=108;	reg signed [w10-1:0] kb310=-82;	reg signed [w10-1:0] kc310=111;	reg signed [w10-1:0] kd310=-76;	reg signed [w10-1:0] ke310=-152;	reg signed [w10-1:0] kf310=-119;	reg signed [w10-1:0] kg310=-68;	reg signed [w10-1:0] kh310=-82;	reg signed [w10-1:0] ki310=44;
reg signed [w10-1:0] ka311=-88;	reg signed [w10-1:0] kb311=-79;	reg signed [w10-1:0] kc311=-144;	reg signed [w10-1:0] kd311=31;	reg signed [w10-1:0] ke311=27;	reg signed [w10-1:0] kf311=-118;	reg signed [w10-1:0] kg311=-31;	reg signed [w10-1:0] kh311=50;	reg signed [w10-1:0] ki311=23;
reg signed [w10-1:0] ka312=-69;	reg signed [w10-1:0] kb312=13;	reg signed [w10-1:0] kc312=101;	reg signed [w10-1:0] kd312=-14;	reg signed [w10-1:0] ke312=24;	reg signed [w10-1:0] kf312=-63;	reg signed [w10-1:0] kg312=64;	reg signed [w10-1:0] kh312=39;	reg signed [w10-1:0] ki312=27;
reg signed [w10-1:0] ka313=11;	reg signed [w10-1:0] kb313=63;	reg signed [w10-1:0] kc313=100;	reg signed [w10-1:0] kd313=15;	reg signed [w10-1:0] ke313=-58;	reg signed [w10-1:0] kf313=-115;	reg signed [w10-1:0] kg313=-108;	reg signed [w10-1:0] kh313=-97;	reg signed [w10-1:0] ki313=-95;
reg signed [w10-1:0] ka314=-34;	reg signed [w10-1:0] kb314=40;	reg signed [w10-1:0] kc314=-11;	reg signed [w10-1:0] kd314=-97;	reg signed [w10-1:0] ke314=43;	reg signed [w10-1:0] kf314=-113;	reg signed [w10-1:0] kg314=115;	reg signed [w10-1:0] kh314=-34;	reg signed [w10-1:0] ki314=-55;
reg signed [w10-1:0] ka315=124;	reg signed [w10-1:0] kb315=51;	reg signed [w10-1:0] kc315=65;	reg signed [w10-1:0] kd315=-114;	reg signed [w10-1:0] ke315=-9;	reg signed [w10-1:0] kf315=-22;	reg signed [w10-1:0] kg315=-94;	reg signed [w10-1:0] kh315=71;	reg signed [w10-1:0] ki315=130;
reg signed [w10-1:0] ka316=-38;	reg signed [w10-1:0] kb316=-34;	reg signed [w10-1:0] kc316=-68;	reg signed [w10-1:0] kd316=93;	reg signed [w10-1:0] ke316=-120;	reg signed [w10-1:0] kf316=-13;	reg signed [w10-1:0] kg316=-18;	reg signed [w10-1:0] kh316=43;	reg signed [w10-1:0] ki316=20;
reg signed [w10-1:0] ka317=-116;	reg signed [w10-1:0] kb317=-43;	reg signed [w10-1:0] kc317=-53;	reg signed [w10-1:0] kd317=111;	reg signed [w10-1:0] ke317=33;	reg signed [w10-1:0] kf317=-22;	reg signed [w10-1:0] kg317=82;	reg signed [w10-1:0] kh317=23;	reg signed [w10-1:0] ki317=-156;
reg signed [w10-1:0] ka318=21;	reg signed [w10-1:0] kb318=-12;	reg signed [w10-1:0] kc318=63;	reg signed [w10-1:0] kd318=110;	reg signed [w10-1:0] ke318=133;	reg signed [w10-1:0] kf318=84;	reg signed [w10-1:0] kg318=47;	reg signed [w10-1:0] kh318=-105;	reg signed [w10-1:0] ki318=75;
reg signed [w10-1:0] ka319=98;	reg signed [w10-1:0] kb319=9;	reg signed [w10-1:0] kc319=-78;	reg signed [w10-1:0] kd319=-63;	reg signed [w10-1:0] ke319=27;	reg signed [w10-1:0] kf319=-52;	reg signed [w10-1:0] kg319=63;	reg signed [w10-1:0] kh319=-14;	reg signed [w10-1:0] ki319=34;
reg signed [w10-1:0] ka320=-35;	reg signed [w10-1:0] kb320=-85;	reg signed [w10-1:0] kc320=-99;	reg signed [w10-1:0] kd320=16;	reg signed [w10-1:0] ke320=42;	reg signed [w10-1:0] kf320=72;	reg signed [w10-1:0] kg320=39;	reg signed [w10-1:0] kh320=62;	reg signed [w10-1:0] ki320=39;
reg signed [w10-1:0] ka321=5;	reg signed [w10-1:0] kb321=-40;	reg signed [w10-1:0] kc321=9;	reg signed [w10-1:0] kd321=35;	reg signed [w10-1:0] ke321=-125;	reg signed [w10-1:0] kf321=-63;	reg signed [w10-1:0] kg321=123;	reg signed [w10-1:0] kh321=36;	reg signed [w10-1:0] ki321=80;
reg signed [w10-1:0] ka322=103;	reg signed [w10-1:0] kb322=14;	reg signed [w10-1:0] kc322=-40;	reg signed [w10-1:0] kd322=8;	reg signed [w10-1:0] ke322=-3;	reg signed [w10-1:0] kf322=91;	reg signed [w10-1:0] kg322=70;	reg signed [w10-1:0] kh322=-121;	reg signed [w10-1:0] ki322=-75;
reg signed [w10-1:0] ka323=-45;	reg signed [w10-1:0] kb323=49;	reg signed [w10-1:0] kc323=108;	reg signed [w10-1:0] kd323=102;	reg signed [w10-1:0] ke323=-70;	reg signed [w10-1:0] kf323=15;	reg signed [w10-1:0] kg323=44;	reg signed [w10-1:0] kh323=-92;	reg signed [w10-1:0] ki323=-145;
reg signed [w10-1:0] ka324=78;	reg signed [w10-1:0] kb324=-84;	reg signed [w10-1:0] kc324=104;	reg signed [w10-1:0] kd324=5;	reg signed [w10-1:0] ke324=31;	reg signed [w10-1:0] kf324=-83;	reg signed [w10-1:0] kg324=176;	reg signed [w10-1:0] kh324=-49;	reg signed [w10-1:0] ki324=60;
reg signed [w10-1:0] ka325=-93;	reg signed [w10-1:0] kb325=-19;	reg signed [w10-1:0] kc325=-44;	reg signed [w10-1:0] kd325=20;	reg signed [w10-1:0] ke325=18;	reg signed [w10-1:0] kf325=59;	reg signed [w10-1:0] kg325=-25;	reg signed [w10-1:0] kh325=-102;	reg signed [w10-1:0] ki325=86;
reg signed [w10-1:0] ka326=-58;	reg signed [w10-1:0] kb326=128;	reg signed [w10-1:0] kc326=42;	reg signed [w10-1:0] kd326=-23;	reg signed [w10-1:0] ke326=75;	reg signed [w10-1:0] kf326=25;	reg signed [w10-1:0] kg326=-104;	reg signed [w10-1:0] kh326=44;	reg signed [w10-1:0] ki326=-24;
reg signed [w10-1:0] ka327=-56;	reg signed [w10-1:0] kb327=83;	reg signed [w10-1:0] kc327=108;	reg signed [w10-1:0] kd327=82;	reg signed [w10-1:0] ke327=-8;	reg signed [w10-1:0] kf327=-46;	reg signed [w10-1:0] kg327=103;	reg signed [w10-1:0] kh327=-27;	reg signed [w10-1:0] ki327=-124;
reg signed [w10-1:0] ka328=-59;	reg signed [w10-1:0] kb328=-38;	reg signed [w10-1:0] kc328=-68;	reg signed [w10-1:0] kd328=-5;	reg signed [w10-1:0] ke328=15;	reg signed [w10-1:0] kf328=30;	reg signed [w10-1:0] kg328=-100;	reg signed [w10-1:0] kh328=-93;	reg signed [w10-1:0] ki328=100;
reg signed [w10-1:0] ka329=68;	reg signed [w10-1:0] kb329=-52;	reg signed [w10-1:0] kc329=58;	reg signed [w10-1:0] kd329=45;	reg signed [w10-1:0] ke329=-65;	reg signed [w10-1:0] kf329=-114;	reg signed [w10-1:0] kg329=74;	reg signed [w10-1:0] kh329=-90;	reg signed [w10-1:0] ki329=-72;
reg signed [w10-1:0] ka330=104;	reg signed [w10-1:0] kb330=-99;	reg signed [w10-1:0] kc330=-7;	reg signed [w10-1:0] kd330=104;	reg signed [w10-1:0] ke330=-59;	reg signed [w10-1:0] kf330=-6;	reg signed [w10-1:0] kg330=108;	reg signed [w10-1:0] kh330=-20;	reg signed [w10-1:0] ki330=28;
reg signed [w10-1:0] ka331=-5;	reg signed [w10-1:0] kb331=17;	reg signed [w10-1:0] kc331=80;	reg signed [w10-1:0] kd331=100;	reg signed [w10-1:0] ke331=-65;	reg signed [w10-1:0] kf331=121;	reg signed [w10-1:0] kg331=45;	reg signed [w10-1:0] kh331=66;	reg signed [w10-1:0] ki331=73;
reg signed [w10-1:0] ka332=-76;	reg signed [w10-1:0] kb332=68;	reg signed [w10-1:0] kc332=-84;	reg signed [w10-1:0] kd332=69;	reg signed [w10-1:0] ke332=-123;	reg signed [w10-1:0] kf332=155;	reg signed [w10-1:0] kg332=-100;	reg signed [w10-1:0] kh332=33;	reg signed [w10-1:0] ki332=-48;
reg signed [w10-1:0] ka333=-91;	reg signed [w10-1:0] kb333=-37;	reg signed [w10-1:0] kc333=-29;	reg signed [w10-1:0] kd333=-25;	reg signed [w10-1:0] ke333=143;	reg signed [w10-1:0] kf333=42;	reg signed [w10-1:0] kg333=34;	reg signed [w10-1:0] kh333=-121;	reg signed [w10-1:0] ki333=-35;
reg signed [w10-1:0] ka334=-122;	reg signed [w10-1:0] kb334=22;	reg signed [w10-1:0] kc334=73;	reg signed [w10-1:0] kd334=42;	reg signed [w10-1:0] ke334=8;	reg signed [w10-1:0] kf334=3;	reg signed [w10-1:0] kg334=-42;	reg signed [w10-1:0] kh334=134;	reg signed [w10-1:0] ki334=-5;
reg signed [w10-1:0] ka335=8;	reg signed [w10-1:0] kb335=-40;	reg signed [w10-1:0] kc335=-77;	reg signed [w10-1:0] kd335=40;	reg signed [w10-1:0] ke335=-22;	reg signed [w10-1:0] kf335=-67;	reg signed [w10-1:0] kg335=-133;	reg signed [w10-1:0] kh335=-70;	reg signed [w10-1:0] ki335=29;
reg signed [w10-1:0] ka336=128;	reg signed [w10-1:0] kb336=-29;	reg signed [w10-1:0] kc336=-42;	reg signed [w10-1:0] kd336=71;	reg signed [w10-1:0] ke336=18;	reg signed [w10-1:0] kf336=82;	reg signed [w10-1:0] kg336=-104;	reg signed [w10-1:0] kh336=-63;	reg signed [w10-1:0] ki336=-73;
reg signed [w10-1:0] ka337=23;	reg signed [w10-1:0] kb337=84;	reg signed [w10-1:0] kc337=130;	reg signed [w10-1:0] kd337=82;	reg signed [w10-1:0] ke337=59;	reg signed [w10-1:0] kf337=28;	reg signed [w10-1:0] kg337=-5;	reg signed [w10-1:0] kh337=-47;	reg signed [w10-1:0] ki337=-71;
reg signed [w10-1:0] ka338=-112;	reg signed [w10-1:0] kb338=-13;	reg signed [w10-1:0] kc338=4;	reg signed [w10-1:0] kd338=-74;	reg signed [w10-1:0] ke338=18;	reg signed [w10-1:0] kf338=5;	reg signed [w10-1:0] kg338=-92;	reg signed [w10-1:0] kh338=133;	reg signed [w10-1:0] ki338=-63;
reg signed [w10-1:0] ka339=-68;	reg signed [w10-1:0] kb339=-19;	reg signed [w10-1:0] kc339=102;	reg signed [w10-1:0] kd339=33;	reg signed [w10-1:0] ke339=-105;	reg signed [w10-1:0] kf339=-17;	reg signed [w10-1:0] kg339=-86;	reg signed [w10-1:0] kh339=-23;	reg signed [w10-1:0] ki339=-93;
reg signed [w10-1:0] ka340=-40;	reg signed [w10-1:0] kb340=-23;	reg signed [w10-1:0] kc340=45;	reg signed [w10-1:0] kd340=33;	reg signed [w10-1:0] ke340=-9;	reg signed [w10-1:0] kf340=45;	reg signed [w10-1:0] kg340=85;	reg signed [w10-1:0] kh340=-7;	reg signed [w10-1:0] ki340=-119;
reg signed [w10-1:0] ka341=126;	reg signed [w10-1:0] kb341=146;	reg signed [w10-1:0] kc341=-32;	reg signed [w10-1:0] kd341=-14;	reg signed [w10-1:0] ke341=139;	reg signed [w10-1:0] kf341=66;	reg signed [w10-1:0] kg341=-29;	reg signed [w10-1:0] kh341=39;	reg signed [w10-1:0] ki341=-9;
reg signed [w10-1:0] ka342=-29;	reg signed [w10-1:0] kb342=-112;	reg signed [w10-1:0] kc342=-119;	reg signed [w10-1:0] kd342=59;	reg signed [w10-1:0] ke342=-35;	reg signed [w10-1:0] kf342=3;	reg signed [w10-1:0] kg342=-39;	reg signed [w10-1:0] kh342=-13;	reg signed [w10-1:0] ki342=109;
reg signed [w10-1:0] ka343=50;	reg signed [w10-1:0] kb343=-139;	reg signed [w10-1:0] kc343=-73;	reg signed [w10-1:0] kd343=-38;	reg signed [w10-1:0] ke343=45;	reg signed [w10-1:0] kf343=33;	reg signed [w10-1:0] kg343=34;	reg signed [w10-1:0] kh343=-26;	reg signed [w10-1:0] ki343=-13;
reg signed [w10-1:0] ka344=-63;	reg signed [w10-1:0] kb344=-94;	reg signed [w10-1:0] kc344=-42;	reg signed [w10-1:0] kd344=0;	reg signed [w10-1:0] ke344=-22;	reg signed [w10-1:0] kf344=-124;	reg signed [w10-1:0] kg344=-77;	reg signed [w10-1:0] kh344=-84;	reg signed [w10-1:0] ki344=-109;
reg signed [w10-1:0] ka345=-58;	reg signed [w10-1:0] kb345=-33;	reg signed [w10-1:0] kc345=-26;	reg signed [w10-1:0] kd345=-44;	reg signed [w10-1:0] ke345=67;	reg signed [w10-1:0] kf345=150;	reg signed [w10-1:0] kg345=31;	reg signed [w10-1:0] kh345=30;	reg signed [w10-1:0] ki345=-56;
reg signed [w10-1:0] ka346=101;	reg signed [w10-1:0] kb346=-107;	reg signed [w10-1:0] kc346=85;	reg signed [w10-1:0] kd346=58;	reg signed [w10-1:0] ke346=-36;	reg signed [w10-1:0] kf346=-59;	reg signed [w10-1:0] kg346=-7;	reg signed [w10-1:0] kh346=144;	reg signed [w10-1:0] ki346=49;
reg signed [w10-1:0] ka347=-140;	reg signed [w10-1:0] kb347=-16;	reg signed [w10-1:0] kc347=48;	reg signed [w10-1:0] kd347=45;	reg signed [w10-1:0] ke347=-100;	reg signed [w10-1:0] kf347=-71;	reg signed [w10-1:0] kg347=88;	reg signed [w10-1:0] kh347=71;	reg signed [w10-1:0] ki347=128;
reg signed [w10-1:0] ka348=-31;	reg signed [w10-1:0] kb348=12;	reg signed [w10-1:0] kc348=-29;	reg signed [w10-1:0] kd348=-2;	reg signed [w10-1:0] ke348=91;	reg signed [w10-1:0] kf348=28;	reg signed [w10-1:0] kg348=-114;	reg signed [w10-1:0] kh348=-17;	reg signed [w10-1:0] ki348=-75;
reg signed [w10-1:0] ka349=19;	reg signed [w10-1:0] kb349=-54;	reg signed [w10-1:0] kc349=-95;	reg signed [w10-1:0] kd349=118;	reg signed [w10-1:0] ke349=82;	reg signed [w10-1:0] kf349=15;	reg signed [w10-1:0] kg349=-5;	reg signed [w10-1:0] kh349=-32;	reg signed [w10-1:0] ki349=-33;
reg signed [w10-1:0] ka350=100;	reg signed [w10-1:0] kb350=8;	reg signed [w10-1:0] kc350=-8;	reg signed [w10-1:0] kd350=47;	reg signed [w10-1:0] ke350=-115;	reg signed [w10-1:0] kf350=77;	reg signed [w10-1:0] kg350=-77;	reg signed [w10-1:0] kh350=-45;	reg signed [w10-1:0] ki350=81;
reg signed [w10-1:0] ka351=-22;	reg signed [w10-1:0] kb351=8;	reg signed [w10-1:0] kc351=-43;	reg signed [w10-1:0] kd351=65;	reg signed [w10-1:0] ke351=16;	reg signed [w10-1:0] kf351=-135;	reg signed [w10-1:0] kg351=-11;	reg signed [w10-1:0] kh351=93;	reg signed [w10-1:0] ki351=-12;
reg signed [w10-1:0] ka352=-48;	reg signed [w10-1:0] kb352=4;	reg signed [w10-1:0] kc352=-49;	reg signed [w10-1:0] kd352=62;	reg signed [w10-1:0] ke352=11;	reg signed [w10-1:0] kf352=23;	reg signed [w10-1:0] kg352=-62;	reg signed [w10-1:0] kh352=-60;	reg signed [w10-1:0] ki352=38;
reg signed [w10-1:0] ka353=-38;	reg signed [w10-1:0] kb353=-48;	reg signed [w10-1:0] kc353=78;	reg signed [w10-1:0] kd353=84;	reg signed [w10-1:0] ke353=-83;	reg signed [w10-1:0] kf353=-50;	reg signed [w10-1:0] kg353=-18;	reg signed [w10-1:0] kh353=23;	reg signed [w10-1:0] ki353=-104;
reg signed [w10-1:0] ka354=29;	reg signed [w10-1:0] kb354=118;	reg signed [w10-1:0] kc354=-56;	reg signed [w10-1:0] kd354=22;	reg signed [w10-1:0] ke354=92;	reg signed [w10-1:0] kf354=93;	reg signed [w10-1:0] kg354=-61;	reg signed [w10-1:0] kh354=-42;	reg signed [w10-1:0] ki354=35;
reg signed [w10-1:0] ka355=150;	reg signed [w10-1:0] kb355=-3;	reg signed [w10-1:0] kc355=63;	reg signed [w10-1:0] kd355=35;	reg signed [w10-1:0] ke355=-135;	reg signed [w10-1:0] kf355=35;	reg signed [w10-1:0] kg355=24;	reg signed [w10-1:0] kh355=-9;	reg signed [w10-1:0] ki355=-83;
reg signed [w10-1:0] ka356=-76;	reg signed [w10-1:0] kb356=-9;	reg signed [w10-1:0] kc356=102;	reg signed [w10-1:0] kd356=34;	reg signed [w10-1:0] ke356=-55;	reg signed [w10-1:0] kf356=-2;	reg signed [w10-1:0] kg356=-17;	reg signed [w10-1:0] kh356=-97;	reg signed [w10-1:0] ki356=-96;
reg signed [w10-1:0] ka357=1;	reg signed [w10-1:0] kb357=-43;	reg signed [w10-1:0] kc357=-52;	reg signed [w10-1:0] kd357=-161;	reg signed [w10-1:0] ke357=36;	reg signed [w10-1:0] kf357=-11;	reg signed [w10-1:0] kg357=20;	reg signed [w10-1:0] kh357=-54;	reg signed [w10-1:0] ki357=-94;
reg signed [w10-1:0] ka358=17;	reg signed [w10-1:0] kb358=84;	reg signed [w10-1:0] kc358=-90;	reg signed [w10-1:0] kd358=64;	reg signed [w10-1:0] ke358=101;	reg signed [w10-1:0] kf358=-39;	reg signed [w10-1:0] kg358=-86;	reg signed [w10-1:0] kh358=36;	reg signed [w10-1:0] ki358=148;
reg signed [w10-1:0] ka359=-31;	reg signed [w10-1:0] kb359=-32;	reg signed [w10-1:0] kc359=127;	reg signed [w10-1:0] kd359=69;	reg signed [w10-1:0] ke359=-37;	reg signed [w10-1:0] kf359=-18;	reg signed [w10-1:0] kg359=-71;	reg signed [w10-1:0] kh359=-4;	reg signed [w10-1:0] ki359=-70;
reg signed [w10-1:0] ka360=-87;	reg signed [w10-1:0] kb360=1;	reg signed [w10-1:0] kc360=34;	reg signed [w10-1:0] kd360=-54;	reg signed [w10-1:0] ke360=80;	reg signed [w10-1:0] kf360=2;	reg signed [w10-1:0] kg360=154;	reg signed [w10-1:0] kh360=98;	reg signed [w10-1:0] ki360=-26;
reg signed [w10-1:0] ka361=53;	reg signed [w10-1:0] kb361=-56;	reg signed [w10-1:0] kc361=-69;	reg signed [w10-1:0] kd361=-56;	reg signed [w10-1:0] ke361=9;	reg signed [w10-1:0] kf361=30;	reg signed [w10-1:0] kg361=36;	reg signed [w10-1:0] kh361=-69;	reg signed [w10-1:0] ki361=109;
reg signed [w10-1:0] ka362=-50;	reg signed [w10-1:0] kb362=85;	reg signed [w10-1:0] kc362=100;	reg signed [w10-1:0] kd362=83;	reg signed [w10-1:0] ke362=63;	reg signed [w10-1:0] kf362=75;	reg signed [w10-1:0] kg362=99;	reg signed [w10-1:0] kh362=-65;	reg signed [w10-1:0] ki362=67;
reg signed [w10-1:0] ka363=88;	reg signed [w10-1:0] kb363=82;	reg signed [w10-1:0] kc363=1;	reg signed [w10-1:0] kd363=0;	reg signed [w10-1:0] ke363=-99;	reg signed [w10-1:0] kf363=9;	reg signed [w10-1:0] kg363=120;	reg signed [w10-1:0] kh363=45;	reg signed [w10-1:0] ki363=81;
reg signed [w10-1:0] ka364=43;	reg signed [w10-1:0] kb364=-82;	reg signed [w10-1:0] kc364=-18;	reg signed [w10-1:0] kd364=112;	reg signed [w10-1:0] ke364=-50;	reg signed [w10-1:0] kf364=-46;	reg signed [w10-1:0] kg364=-46;	reg signed [w10-1:0] kh364=-39;	reg signed [w10-1:0] ki364=77;
reg signed [w10-1:0] ka365=59;	reg signed [w10-1:0] kb365=-96;	reg signed [w10-1:0] kc365=-4;	reg signed [w10-1:0] kd365=75;	reg signed [w10-1:0] ke365=-104;	reg signed [w10-1:0] kf365=-40;	reg signed [w10-1:0] kg365=-79;	reg signed [w10-1:0] kh365=37;	reg signed [w10-1:0] ki365=-134;
reg signed [w10-1:0] ka366=-81;	reg signed [w10-1:0] kb366=57;	reg signed [w10-1:0] kc366=-59;	reg signed [w10-1:0] kd366=37;	reg signed [w10-1:0] ke366=151;	reg signed [w10-1:0] kf366=-34;	reg signed [w10-1:0] kg366=75;	reg signed [w10-1:0] kh366=45;	reg signed [w10-1:0] ki366=-91;
reg signed [w10-1:0] ka367=26;	reg signed [w10-1:0] kb367=93;	reg signed [w10-1:0] kc367=-98;	reg signed [w10-1:0] kd367=-96;	reg signed [w10-1:0] ke367=-5;	reg signed [w10-1:0] kf367=-61;	reg signed [w10-1:0] kg367=-105;	reg signed [w10-1:0] kh367=56;	reg signed [w10-1:0] ki367=-4;
reg signed [w10-1:0] ka368=83;	reg signed [w10-1:0] kb368=-32;	reg signed [w10-1:0] kc368=-76;	reg signed [w10-1:0] kd368=109;	reg signed [w10-1:0] ke368=-108;	reg signed [w10-1:0] kf368=70;	reg signed [w10-1:0] kg368=-15;	reg signed [w10-1:0] kh368=81;	reg signed [w10-1:0] ki368=-48;
reg signed [w10-1:0] ka369=-8;	reg signed [w10-1:0] kb369=71;	reg signed [w10-1:0] kc369=53;	reg signed [w10-1:0] kd369=-73;	reg signed [w10-1:0] ke369=99;	reg signed [w10-1:0] kf369=17;	reg signed [w10-1:0] kg369=-96;	reg signed [w10-1:0] kh369=-10;	reg signed [w10-1:0] ki369=-103;
reg signed [w10-1:0] ka370=-111;	reg signed [w10-1:0] kb370=54;	reg signed [w10-1:0] kc370=56;	reg signed [w10-1:0] kd370=-73;	reg signed [w10-1:0] ke370=91;	reg signed [w10-1:0] kf370=-76;	reg signed [w10-1:0] kg370=-36;	reg signed [w10-1:0] kh370=-130;	reg signed [w10-1:0] ki370=35;
reg signed [w10-1:0] ka371=-114;	reg signed [w10-1:0] kb371=5;	reg signed [w10-1:0] kc371=25;	reg signed [w10-1:0] kd371=-40;	reg signed [w10-1:0] ke371=103;	reg signed [w10-1:0] kf371=-73;	reg signed [w10-1:0] kg371=56;	reg signed [w10-1:0] kh371=-58;	reg signed [w10-1:0] ki371=-37;
reg signed [w10-1:0] ka372=98;	reg signed [w10-1:0] kb372=64;	reg signed [w10-1:0] kc372=36;	reg signed [w10-1:0] kd372=-33;	reg signed [w10-1:0] ke372=-102;	reg signed [w10-1:0] kf372=-34;	reg signed [w10-1:0] kg372=100;	reg signed [w10-1:0] kh372=-26;	reg signed [w10-1:0] ki372=-80;
reg signed [w10-1:0] ka373=-18;	reg signed [w10-1:0] kb373=117;	reg signed [w10-1:0] kc373=86;	reg signed [w10-1:0] kd373=75;	reg signed [w10-1:0] ke373=59;	reg signed [w10-1:0] kf373=50;	reg signed [w10-1:0] kg373=93;	reg signed [w10-1:0] kh373=34;	reg signed [w10-1:0] ki373=31;
reg signed [w10-1:0] ka374=-92;	reg signed [w10-1:0] kb374=-77;	reg signed [w10-1:0] kc374=-57;	reg signed [w10-1:0] kd374=-96;	reg signed [w10-1:0] ke374=-24;	reg signed [w10-1:0] kf374=111;	reg signed [w10-1:0] kg374=9;	reg signed [w10-1:0] kh374=-72;	reg signed [w10-1:0] ki374=72;
reg signed [w10-1:0] ka375=117;	reg signed [w10-1:0] kb375=97;	reg signed [w10-1:0] kc375=-58;	reg signed [w10-1:0] kd375=-82;	reg signed [w10-1:0] ke375=57;	reg signed [w10-1:0] kf375=4;	reg signed [w10-1:0] kg375=-110;	reg signed [w10-1:0] kh375=8;	reg signed [w10-1:0] ki375=-123;
reg signed [w10-1:0] ka376=-1;	reg signed [w10-1:0] kb376=140;	reg signed [w10-1:0] kc376=-36;	reg signed [w10-1:0] kd376=-119;	reg signed [w10-1:0] ke376=63;	reg signed [w10-1:0] kf376=47;	reg signed [w10-1:0] kg376=-41;	reg signed [w10-1:0] kh376=-27;	reg signed [w10-1:0] ki376=39;
reg signed [w10-1:0] ka377=-102;	reg signed [w10-1:0] kb377=52;	reg signed [w10-1:0] kc377=34;	reg signed [w10-1:0] kd377=-48;	reg signed [w10-1:0] ke377=87;	reg signed [w10-1:0] kf377=-89;	reg signed [w10-1:0] kg377=-108;	reg signed [w10-1:0] kh377=-53;	reg signed [w10-1:0] ki377=-37;
reg signed [w10-1:0] ka378=53;	reg signed [w10-1:0] kb378=87;	reg signed [w10-1:0] kc378=-37;	reg signed [w10-1:0] kd378=35;	reg signed [w10-1:0] ke378=-53;	reg signed [w10-1:0] kf378=85;	reg signed [w10-1:0] kg378=52;	reg signed [w10-1:0] kh378=26;	reg signed [w10-1:0] ki378=41;
reg signed [w10-1:0] ka379=73;	reg signed [w10-1:0] kb379=-14;	reg signed [w10-1:0] kc379=76;	reg signed [w10-1:0] kd379=53;	reg signed [w10-1:0] ke379=-94;	reg signed [w10-1:0] kf379=-132;	reg signed [w10-1:0] kg379=62;	reg signed [w10-1:0] kh379=-96;	reg signed [w10-1:0] ki379=-10;
reg signed [w10-1:0] ka380=56;	reg signed [w10-1:0] kb380=-124;	reg signed [w10-1:0] kc380=-54;	reg signed [w10-1:0] kd380=122;	reg signed [w10-1:0] ke380=-11;	reg signed [w10-1:0] kf380=123;	reg signed [w10-1:0] kg380=2;	reg signed [w10-1:0] kh380=-100;	reg signed [w10-1:0] ki380=-73;
reg signed [w10-1:0] ka381=57;	reg signed [w10-1:0] kb381=-95;	reg signed [w10-1:0] kc381=-87;	reg signed [w10-1:0] kd381=-67;	reg signed [w10-1:0] ke381=-114;	reg signed [w10-1:0] kf381=71;	reg signed [w10-1:0] kg381=1;	reg signed [w10-1:0] kh381=92;	reg signed [w10-1:0] ki381=-55;
reg signed [w10-1:0] ka382=-12;	reg signed [w10-1:0] kb382=66;	reg signed [w10-1:0] kc382=93;	reg signed [w10-1:0] kd382=-46;	reg signed [w10-1:0] ke382=-22;	reg signed [w10-1:0] kf382=33;	reg signed [w10-1:0] kg382=-135;	reg signed [w10-1:0] kh382=24;	reg signed [w10-1:0] ki382=-43;
reg signed [w10-1:0] ka383=41;	reg signed [w10-1:0] kb383=-6;	reg signed [w10-1:0] kc383=-118;	reg signed [w10-1:0] kd383=-118;	reg signed [w10-1:0] ke383=-101;	reg signed [w10-1:0] kf383=-98;	reg signed [w10-1:0] kg383=-87;	reg signed [w10-1:0] kh383=94;	reg signed [w10-1:0] ki383=-9;
reg signed [w10-1:0] ka384=-65;	reg signed [w10-1:0] kb384=-18;	reg signed [w10-1:0] kc384=12;	reg signed [w10-1:0] kd384=127;	reg signed [w10-1:0] ke384=-71;	reg signed [w10-1:0] kf384=107;	reg signed [w10-1:0] kg384=-22;	reg signed [w10-1:0] kh384=-6;	reg signed [w10-1:0] ki384=5;
reg signed [w10-1:0] ka385=90;	reg signed [w10-1:0] kb385=-96;	reg signed [w10-1:0] kc385=58;	reg signed [w10-1:0] kd385=-109;	reg signed [w10-1:0] ke385=25;	reg signed [w10-1:0] kf385=-103;	reg signed [w10-1:0] kg385=-42;	reg signed [w10-1:0] kh385=36;	reg signed [w10-1:0] ki385=10;
reg signed [w10-1:0] ka386=-33;	reg signed [w10-1:0] kb386=-84;	reg signed [w10-1:0] kc386=39;	reg signed [w10-1:0] kd386=-31;	reg signed [w10-1:0] ke386=-64;	reg signed [w10-1:0] kf386=-51;	reg signed [w10-1:0] kg386=29;	reg signed [w10-1:0] kh386=-31;	reg signed [w10-1:0] ki386=-37;
reg signed [w10-1:0] ka387=-23;	reg signed [w10-1:0] kb387=-66;	reg signed [w10-1:0] kc387=71;	reg signed [w10-1:0] kd387=94;	reg signed [w10-1:0] ke387=41;	reg signed [w10-1:0] kf387=-104;	reg signed [w10-1:0] kg387=44;	reg signed [w10-1:0] kh387=-102;	reg signed [w10-1:0] ki387=-3;
reg signed [w10-1:0] ka388=27;	reg signed [w10-1:0] kb388=-86;	reg signed [w10-1:0] kc388=-39;	reg signed [w10-1:0] kd388=-132;	reg signed [w10-1:0] ke388=11;	reg signed [w10-1:0] kf388=76;	reg signed [w10-1:0] kg388=15;	reg signed [w10-1:0] kh388=-49;	reg signed [w10-1:0] ki388=-106;
reg signed [w10-1:0] ka389=49;	reg signed [w10-1:0] kb389=-45;	reg signed [w10-1:0] kc389=68;	reg signed [w10-1:0] kd389=-58;	reg signed [w10-1:0] ke389=-33;	reg signed [w10-1:0] kf389=92;	reg signed [w10-1:0] kg389=136;	reg signed [w10-1:0] kh389=150;	reg signed [w10-1:0] ki389=121;
reg signed [w10-1:0] ka390=-94;	reg signed [w10-1:0] kb390=26;	reg signed [w10-1:0] kc390=-5;	reg signed [w10-1:0] kd390=-18;	reg signed [w10-1:0] ke390=85;	reg signed [w10-1:0] kf390=-92;	reg signed [w10-1:0] kg390=34;	reg signed [w10-1:0] kh390=-66;	reg signed [w10-1:0] ki390=-126;
reg signed [w10-1:0] ka391=75;	reg signed [w10-1:0] kb391=-37;	reg signed [w10-1:0] kc391=28;	reg signed [w10-1:0] kd391=-69;	reg signed [w10-1:0] ke391=-77;	reg signed [w10-1:0] kf391=-104;	reg signed [w10-1:0] kg391=-117;	reg signed [w10-1:0] kh391=-107;	reg signed [w10-1:0] ki391=99;
reg signed [w10-1:0] ka392=-115;	reg signed [w10-1:0] kb392=-13;	reg signed [w10-1:0] kc392=113;	reg signed [w10-1:0] kd392=6;	reg signed [w10-1:0] ke392=74;	reg signed [w10-1:0] kf392=-34;	reg signed [w10-1:0] kg392=-83;	reg signed [w10-1:0] kh392=29;	reg signed [w10-1:0] ki392=-46;
reg signed [w10-1:0] ka393=31;	reg signed [w10-1:0] kb393=-69;	reg signed [w10-1:0] kc393=-46;	reg signed [w10-1:0] kd393=50;	reg signed [w10-1:0] ke393=-87;	reg signed [w10-1:0] kf393=-97;	reg signed [w10-1:0] kg393=-17;	reg signed [w10-1:0] kh393=-90;	reg signed [w10-1:0] ki393=-115;
reg signed [w10-1:0] ka394=144;	reg signed [w10-1:0] kb394=85;	reg signed [w10-1:0] kc394=74;	reg signed [w10-1:0] kd394=132;	reg signed [w10-1:0] ke394=-37;	reg signed [w10-1:0] kf394=-5;	reg signed [w10-1:0] kg394=4;	reg signed [w10-1:0] kh394=15;	reg signed [w10-1:0] ki394=2;
reg signed [w10-1:0] ka395=-98;	reg signed [w10-1:0] kb395=61;	reg signed [w10-1:0] kc395=-70;	reg signed [w10-1:0] kd395=64;	reg signed [w10-1:0] ke395=-68;	reg signed [w10-1:0] kf395=-52;	reg signed [w10-1:0] kg395=38;	reg signed [w10-1:0] kh395=92;	reg signed [w10-1:0] ki395=-53;
reg signed [w10-1:0] ka396=-7;	reg signed [w10-1:0] kb396=-129;	reg signed [w10-1:0] kc396=-74;	reg signed [w10-1:0] kd396=-84;	reg signed [w10-1:0] ke396=-5;	reg signed [w10-1:0] kf396=-128;	reg signed [w10-1:0] kg396=82;	reg signed [w10-1:0] kh396=3;	reg signed [w10-1:0] ki396=74;
reg signed [w10-1:0] ka397=83;	reg signed [w10-1:0] kb397=17;	reg signed [w10-1:0] kc397=122;	reg signed [w10-1:0] kd397=-43;	reg signed [w10-1:0] ke397=98;	reg signed [w10-1:0] kf397=90;	reg signed [w10-1:0] kg397=-45;	reg signed [w10-1:0] kh397=67;	reg signed [w10-1:0] ki397=3;
reg signed [w10-1:0] ka398=107;	reg signed [w10-1:0] kb398=0;	reg signed [w10-1:0] kc398=-60;	reg signed [w10-1:0] kd398=-30;	reg signed [w10-1:0] ke398=95;	reg signed [w10-1:0] kf398=137;	reg signed [w10-1:0] kg398=95;	reg signed [w10-1:0] kh398=36;	reg signed [w10-1:0] ki398=26;
reg signed [w10-1:0] ka399=54;	reg signed [w10-1:0] kb399=-89;	reg signed [w10-1:0] kc399=-17;	reg signed [w10-1:0] kd399=2;	reg signed [w10-1:0] ke399=75;	reg signed [w10-1:0] kf399=59;	reg signed [w10-1:0] kg399=110;	reg signed [w10-1:0] kh399=-97;	reg signed [w10-1:0] ki399=-43;
reg signed [w10-1:0] ka400=56;	reg signed [w10-1:0] kb400=24;	reg signed [w10-1:0] kc400=51;	reg signed [w10-1:0] kd400=-124;	reg signed [w10-1:0] ke400=86;	reg signed [w10-1:0] kf400=48;	reg signed [w10-1:0] kg400=-103;	reg signed [w10-1:0] kh400=-69;	reg signed [w10-1:0] ki400=12;
reg signed [w10-1:0] ka401=-99;	reg signed [w10-1:0] kb401=30;	reg signed [w10-1:0] kc401=-10;	reg signed [w10-1:0] kd401=-59;	reg signed [w10-1:0] ke401=49;	reg signed [w10-1:0] kf401=87;	reg signed [w10-1:0] kg401=-68;	reg signed [w10-1:0] kh401=114;	reg signed [w10-1:0] ki401=84;
reg signed [w10-1:0] ka402=-96;	reg signed [w10-1:0] kb402=-107;	reg signed [w10-1:0] kc402=15;	reg signed [w10-1:0] kd402=-50;	reg signed [w10-1:0] ke402=-30;	reg signed [w10-1:0] kf402=12;	reg signed [w10-1:0] kg402=-37;	reg signed [w10-1:0] kh402=-20;	reg signed [w10-1:0] ki402=15;
reg signed [w10-1:0] ka403=-31;	reg signed [w10-1:0] kb403=19;	reg signed [w10-1:0] kc403=-6;	reg signed [w10-1:0] kd403=66;	reg signed [w10-1:0] ke403=60;	reg signed [w10-1:0] kf403=54;	reg signed [w10-1:0] kg403=-100;	reg signed [w10-1:0] kh403=-54;	reg signed [w10-1:0] ki403=10;
reg signed [w10-1:0] ka404=72;	reg signed [w10-1:0] kb404=-20;	reg signed [w10-1:0] kc404=-26;	reg signed [w10-1:0] kd404=34;	reg signed [w10-1:0] ke404=-132;	reg signed [w10-1:0] kf404=-24;	reg signed [w10-1:0] kg404=149;	reg signed [w10-1:0] kh404=118;	reg signed [w10-1:0] ki404=33;
reg signed [w10-1:0] ka405=-174;	reg signed [w10-1:0] kb405=-191;	reg signed [w10-1:0] kc405=-60;	reg signed [w10-1:0] kd405=-132;	reg signed [w10-1:0] ke405=-168;	reg signed [w10-1:0] kf405=10;	reg signed [w10-1:0] kg405=47;	reg signed [w10-1:0] kh405=-108;	reg signed [w10-1:0] ki405=-136;
reg signed [w10-1:0] ka406=-55;	reg signed [w10-1:0] kb406=-61;	reg signed [w10-1:0] kc406=26;	reg signed [w10-1:0] kd406=57;	reg signed [w10-1:0] ke406=102;	reg signed [w10-1:0] kf406=127;	reg signed [w10-1:0] kg406=64;	reg signed [w10-1:0] kh406=70;	reg signed [w10-1:0] ki406=5;
reg signed [w10-1:0] ka407=-61;	reg signed [w10-1:0] kb407=-43;	reg signed [w10-1:0] kc407=-86;	reg signed [w10-1:0] kd407=114;	reg signed [w10-1:0] ke407=19;	reg signed [w10-1:0] kf407=-10;	reg signed [w10-1:0] kg407=88;	reg signed [w10-1:0] kh407=-62;	reg signed [w10-1:0] ki407=5;
reg signed [w10-1:0] ka408=-16;	reg signed [w10-1:0] kb408=97;	reg signed [w10-1:0] kc408=-4;	reg signed [w10-1:0] kd408=-27;	reg signed [w10-1:0] ke408=68;	reg signed [w10-1:0] kf408=-91;	reg signed [w10-1:0] kg408=-106;	reg signed [w10-1:0] kh408=-60;	reg signed [w10-1:0] ki408=-75;
reg signed [w10-1:0] ka409=62;	reg signed [w10-1:0] kb409=63;	reg signed [w10-1:0] kc409=-39;	reg signed [w10-1:0] kd409=-99;	reg signed [w10-1:0] ke409=7;	reg signed [w10-1:0] kf409=-47;	reg signed [w10-1:0] kg409=-61;	reg signed [w10-1:0] kh409=9;	reg signed [w10-1:0] ki409=-28;
reg signed [w10-1:0] ka410=12;	reg signed [w10-1:0] kb410=-9;	reg signed [w10-1:0] kc410=-69;	reg signed [w10-1:0] kd410=69;	reg signed [w10-1:0] ke410=121;	reg signed [w10-1:0] kf410=-53;	reg signed [w10-1:0] kg410=22;	reg signed [w10-1:0] kh410=-18;	reg signed [w10-1:0] ki410=-95;
reg signed [w10-1:0] ka411=-31;	reg signed [w10-1:0] kb411=-56;	reg signed [w10-1:0] kc411=-73;	reg signed [w10-1:0] kd411=15;	reg signed [w10-1:0] ke411=-67;	reg signed [w10-1:0] kf411=-69;	reg signed [w10-1:0] kg411=70;	reg signed [w10-1:0] kh411=25;	reg signed [w10-1:0] ki411=-161;
reg signed [w10-1:0] ka412=5;	reg signed [w10-1:0] kb412=55;	reg signed [w10-1:0] kc412=119;	reg signed [w10-1:0] kd412=-98;	reg signed [w10-1:0] ke412=-43;	reg signed [w10-1:0] kf412=57;	reg signed [w10-1:0] kg412=-51;	reg signed [w10-1:0] kh412=-2;	reg signed [w10-1:0] ki412=-1;
reg signed [w10-1:0] ka413=0;	reg signed [w10-1:0] kb413=42;	reg signed [w10-1:0] kc413=50;	reg signed [w10-1:0] kd413=-35;	reg signed [w10-1:0] ke413=118;	reg signed [w10-1:0] kf413=43;	reg signed [w10-1:0] kg413=-111;	reg signed [w10-1:0] kh413=69;	reg signed [w10-1:0] ki413=30;
reg signed [w10-1:0] ka414=-46;	reg signed [w10-1:0] kb414=46;	reg signed [w10-1:0] kc414=116;	reg signed [w10-1:0] kd414=48;	reg signed [w10-1:0] ke414=-91;	reg signed [w10-1:0] kf414=73;	reg signed [w10-1:0] kg414=-9;	reg signed [w10-1:0] kh414=-120;	reg signed [w10-1:0] ki414=55;
reg signed [w10-1:0] ka415=-80;	reg signed [w10-1:0] kb415=92;	reg signed [w10-1:0] kc415=37;	reg signed [w10-1:0] kd415=-8;	reg signed [w10-1:0] ke415=82;	reg signed [w10-1:0] kf415=-131;	reg signed [w10-1:0] kg415=166;	reg signed [w10-1:0] kh415=-22;	reg signed [w10-1:0] ki415=40;
reg signed [w10-1:0] ka416=11;	reg signed [w10-1:0] kb416=-90;	reg signed [w10-1:0] kc416=-89;	reg signed [w10-1:0] kd416=60;	reg signed [w10-1:0] ke416=-14;	reg signed [w10-1:0] kf416=34;	reg signed [w10-1:0] kg416=-4;	reg signed [w10-1:0] kh416=-64;	reg signed [w10-1:0] ki416=-127;
reg signed [w10-1:0] ka417=102;	reg signed [w10-1:0] kb417=-20;	reg signed [w10-1:0] kc417=76;	reg signed [w10-1:0] kd417=113;	reg signed [w10-1:0] ke417=-64;	reg signed [w10-1:0] kf417=37;	reg signed [w10-1:0] kg417=-59;	reg signed [w10-1:0] kh417=78;	reg signed [w10-1:0] ki417=-44;
reg signed [w10-1:0] ka418=20;	reg signed [w10-1:0] kb418=107;	reg signed [w10-1:0] kc418=-47;	reg signed [w10-1:0] kd418=-19;	reg signed [w10-1:0] ke418=-44;	reg signed [w10-1:0] kf418=-16;	reg signed [w10-1:0] kg418=68;	reg signed [w10-1:0] kh418=54;	reg signed [w10-1:0] ki418=89;
reg signed [w10-1:0] ka419=-14;	reg signed [w10-1:0] kb419=60;	reg signed [w10-1:0] kc419=-48;	reg signed [w10-1:0] kd419=-105;	reg signed [w10-1:0] ke419=47;	reg signed [w10-1:0] kf419=3;	reg signed [w10-1:0] kg419=51;	reg signed [w10-1:0] kh419=105;	reg signed [w10-1:0] ki419=8;
reg signed [w10-1:0] ka420=59;	reg signed [w10-1:0] kb420=-15;	reg signed [w10-1:0] kc420=90;	reg signed [w10-1:0] kd420=-11;	reg signed [w10-1:0] ke420=148;	reg signed [w10-1:0] kf420=115;	reg signed [w10-1:0] kg420=50;	reg signed [w10-1:0] kh420=-4;	reg signed [w10-1:0] ki420=3;
reg signed [w10-1:0] ka421=36;	reg signed [w10-1:0] kb421=-93;	reg signed [w10-1:0] kc421=123;	reg signed [w10-1:0] kd421=98;	reg signed [w10-1:0] ke421=-87;	reg signed [w10-1:0] kf421=20;	reg signed [w10-1:0] kg421=78;	reg signed [w10-1:0] kh421=106;	reg signed [w10-1:0] ki421=130;
reg signed [w10-1:0] ka422=26;	reg signed [w10-1:0] kb422=7;	reg signed [w10-1:0] kc422=-47;	reg signed [w10-1:0] kd422=-14;	reg signed [w10-1:0] ke422=30;	reg signed [w10-1:0] kf422=53;	reg signed [w10-1:0] kg422=-171;	reg signed [w10-1:0] kh422=35;	reg signed [w10-1:0] ki422=-2;
reg signed [w10-1:0] ka423=110;	reg signed [w10-1:0] kb423=-77;	reg signed [w10-1:0] kc423=-116;	reg signed [w10-1:0] kd423=-8;	reg signed [w10-1:0] ke423=-53;	reg signed [w10-1:0] kf423=-110;	reg signed [w10-1:0] kg423=-127;	reg signed [w10-1:0] kh423=-15;	reg signed [w10-1:0] ki423=-29;
reg signed [w10-1:0] ka424=76;	reg signed [w10-1:0] kb424=-73;	reg signed [w10-1:0] kc424=54;	reg signed [w10-1:0] kd424=84;	reg signed [w10-1:0] ke424=-56;	reg signed [w10-1:0] kf424=-78;	reg signed [w10-1:0] kg424=-16;	reg signed [w10-1:0] kh424=-134;	reg signed [w10-1:0] ki424=69;
reg signed [w10-1:0] ka425=-90;	reg signed [w10-1:0] kb425=49;	reg signed [w10-1:0] kc425=46;	reg signed [w10-1:0] kd425=-21;	reg signed [w10-1:0] ke425=52;	reg signed [w10-1:0] kf425=-57;	reg signed [w10-1:0] kg425=-77;	reg signed [w10-1:0] kh425=-58;	reg signed [w10-1:0] ki425=-139;
reg signed [w10-1:0] ka426=85;	reg signed [w10-1:0] kb426=-100;	reg signed [w10-1:0] kc426=25;	reg signed [w10-1:0] kd426=137;	reg signed [w10-1:0] ke426=89;	reg signed [w10-1:0] kf426=-19;	reg signed [w10-1:0] kg426=55;	reg signed [w10-1:0] kh426=120;	reg signed [w10-1:0] ki426=-95;
reg signed [w10-1:0] ka427=1;	reg signed [w10-1:0] kb427=34;	reg signed [w10-1:0] kc427=-88;	reg signed [w10-1:0] kd427=96;	reg signed [w10-1:0] ke427=93;	reg signed [w10-1:0] kf427=-88;	reg signed [w10-1:0] kg427=36;	reg signed [w10-1:0] kh427=-104;	reg signed [w10-1:0] ki427=-128;
reg signed [w10-1:0] ka428=-104;	reg signed [w10-1:0] kb428=29;	reg signed [w10-1:0] kc428=-52;	reg signed [w10-1:0] kd428=53;	reg signed [w10-1:0] ke428=-136;	reg signed [w10-1:0] kf428=7;	reg signed [w10-1:0] kg428=-78;	reg signed [w10-1:0] kh428=1;	reg signed [w10-1:0] ki428=46;
reg signed [w10-1:0] ka429=-75;	reg signed [w10-1:0] kb429=-47;	reg signed [w10-1:0] kc429=47;	reg signed [w10-1:0] kd429=-64;	reg signed [w10-1:0] ke429=54;	reg signed [w10-1:0] kf429=51;	reg signed [w10-1:0] kg429=-85;	reg signed [w10-1:0] kh429=80;	reg signed [w10-1:0] ki429=67;
reg signed [w10-1:0] ka430=-148;	reg signed [w10-1:0] kb430=-128;	reg signed [w10-1:0] kc430=17;	reg signed [w10-1:0] kd430=101;	reg signed [w10-1:0] ke430=-18;	reg signed [w10-1:0] kf430=123;	reg signed [w10-1:0] kg430=28;	reg signed [w10-1:0] kh430=3;	reg signed [w10-1:0] ki430=42;
reg signed [w10-1:0] ka431=50;	reg signed [w10-1:0] kb431=28;	reg signed [w10-1:0] kc431=80;	reg signed [w10-1:0] kd431=80;	reg signed [w10-1:0] ke431=-104;	reg signed [w10-1:0] kf431=-73;	reg signed [w10-1:0] kg431=-81;	reg signed [w10-1:0] kh431=6;	reg signed [w10-1:0] ki431=4;
reg signed [w10-1:0] ka432=-60;	reg signed [w10-1:0] kb432=-99;	reg signed [w10-1:0] kc432=-56;	reg signed [w10-1:0] kd432=50;	reg signed [w10-1:0] ke432=100;	reg signed [w10-1:0] kf432=-113;	reg signed [w10-1:0] kg432=53;	reg signed [w10-1:0] kh432=145;	reg signed [w10-1:0] ki432=128;
reg signed [w10-1:0] ka433=12;	reg signed [w10-1:0] kb433=102;	reg signed [w10-1:0] kc433=68;	reg signed [w10-1:0] kd433=44;	reg signed [w10-1:0] ke433=114;	reg signed [w10-1:0] kf433=156;	reg signed [w10-1:0] kg433=104;	reg signed [w10-1:0] kh433=-27;	reg signed [w10-1:0] ki433=111;
reg signed [w10-1:0] ka434=27;	reg signed [w10-1:0] kb434=-51;	reg signed [w10-1:0] kc434=-35;	reg signed [w10-1:0] kd434=-116;	reg signed [w10-1:0] ke434=-40;	reg signed [w10-1:0] kf434=88;	reg signed [w10-1:0] kg434=61;	reg signed [w10-1:0] kh434=25;	reg signed [w10-1:0] ki434=-73;
reg signed [w10-1:0] ka435=-7;	reg signed [w10-1:0] kb435=-107;	reg signed [w10-1:0] kc435=31;	reg signed [w10-1:0] kd435=-21;	reg signed [w10-1:0] ke435=103;	reg signed [w10-1:0] kf435=-90;	reg signed [w10-1:0] kg435=-12;	reg signed [w10-1:0] kh435=79;	reg signed [w10-1:0] ki435=-7;
reg signed [w10-1:0] ka436=-63;	reg signed [w10-1:0] kb436=62;	reg signed [w10-1:0] kc436=33;	reg signed [w10-1:0] kd436=-141;	reg signed [w10-1:0] ke436=68;	reg signed [w10-1:0] kf436=82;	reg signed [w10-1:0] kg436=-51;	reg signed [w10-1:0] kh436=-109;	reg signed [w10-1:0] ki436=-30;
reg signed [w10-1:0] ka437=-41;	reg signed [w10-1:0] kb437=45;	reg signed [w10-1:0] kc437=-21;	reg signed [w10-1:0] kd437=-210;	reg signed [w10-1:0] ke437=-2;	reg signed [w10-1:0] kf437=-28;	reg signed [w10-1:0] kg437=4;	reg signed [w10-1:0] kh437=-29;	reg signed [w10-1:0] ki437=-83;
reg signed [w10-1:0] ka438=9;	reg signed [w10-1:0] kb438=78;	reg signed [w10-1:0] kc438=68;	reg signed [w10-1:0] kd438=41;	reg signed [w10-1:0] ke438=28;	reg signed [w10-1:0] kf438=-49;	reg signed [w10-1:0] kg438=46;	reg signed [w10-1:0] kh438=48;	reg signed [w10-1:0] ki438=-83;
reg signed [w10-1:0] ka439=-18;	reg signed [w10-1:0] kb439=-96;	reg signed [w10-1:0] kc439=67;	reg signed [w10-1:0] kd439=44;	reg signed [w10-1:0] ke439=-26;	reg signed [w10-1:0] kf439=68;	reg signed [w10-1:0] kg439=-53;	reg signed [w10-1:0] kh439=-75;	reg signed [w10-1:0] ki439=-64;
reg signed [w10-1:0] ka440=102;	reg signed [w10-1:0] kb440=-67;	reg signed [w10-1:0] kc440=22;	reg signed [w10-1:0] kd440=-7;	reg signed [w10-1:0] ke440=-35;	reg signed [w10-1:0] kf440=-88;	reg signed [w10-1:0] kg440=-37;	reg signed [w10-1:0] kh440=73;	reg signed [w10-1:0] ki440=-38;
reg signed [w10-1:0] ka441=-4;	reg signed [w10-1:0] kb441=32;	reg signed [w10-1:0] kc441=-6;	reg signed [w10-1:0] kd441=116;	reg signed [w10-1:0] ke441=52;	reg signed [w10-1:0] kf441=121;	reg signed [w10-1:0] kg441=15;	reg signed [w10-1:0] kh441=-33;	reg signed [w10-1:0] ki441=-103;
reg signed [w10-1:0] ka442=-103;	reg signed [w10-1:0] kb442=7;	reg signed [w10-1:0] kc442=32;	reg signed [w10-1:0] kd442=-40;	reg signed [w10-1:0] ke442=-23;	reg signed [w10-1:0] kf442=40;	reg signed [w10-1:0] kg442=104;	reg signed [w10-1:0] kh442=10;	reg signed [w10-1:0] ki442=86;
reg signed [w10-1:0] ka443=-142;	reg signed [w10-1:0] kb443=-13;	reg signed [w10-1:0] kc443=-41;	reg signed [w10-1:0] kd443=-52;	reg signed [w10-1:0] ke443=-8;	reg signed [w10-1:0] kf443=19;	reg signed [w10-1:0] kg443=56;	reg signed [w10-1:0] kh443=-68;	reg signed [w10-1:0] ki443=28;
reg signed [w10-1:0] ka444=-80;	reg signed [w10-1:0] kb444=78;	reg signed [w10-1:0] kc444=35;	reg signed [w10-1:0] kd444=160;	reg signed [w10-1:0] ke444=15;	reg signed [w10-1:0] kf444=13;	reg signed [w10-1:0] kg444=88;	reg signed [w10-1:0] kh444=-72;	reg signed [w10-1:0] ki444=76;
reg signed [w10-1:0] ka445=33;	reg signed [w10-1:0] kb445=-61;	reg signed [w10-1:0] kc445=-55;	reg signed [w10-1:0] kd445=-107;	reg signed [w10-1:0] ke445=-72;	reg signed [w10-1:0] kf445=-24;	reg signed [w10-1:0] kg445=52;	reg signed [w10-1:0] kh445=-43;	reg signed [w10-1:0] ki445=-74;
reg signed [w10-1:0] ka446=87;	reg signed [w10-1:0] kb446=-13;	reg signed [w10-1:0] kc446=-126;	reg signed [w10-1:0] kd446=-27;	reg signed [w10-1:0] ke446=-96;	reg signed [w10-1:0] kf446=-65;	reg signed [w10-1:0] kg446=-109;	reg signed [w10-1:0] kh446=90;	reg signed [w10-1:0] ki446=-33;
reg signed [w10-1:0] ka447=30;	reg signed [w10-1:0] kb447=-39;	reg signed [w10-1:0] kc447=33;	reg signed [w10-1:0] kd447=-1;	reg signed [w10-1:0] ke447=105;	reg signed [w10-1:0] kf447=-25;	reg signed [w10-1:0] kg447=90;	reg signed [w10-1:0] kh447=-24;	reg signed [w10-1:0] ki447=120;
reg signed [w10-1:0] ka448=-69;	reg signed [w10-1:0] kb448=123;	reg signed [w10-1:0] kc448=28;	reg signed [w10-1:0] kd448=-54;	reg signed [w10-1:0] ke448=-50;	reg signed [w10-1:0] kf448=53;	reg signed [w10-1:0] kg448=-24;	reg signed [w10-1:0] kh448=-32;	reg signed [w10-1:0] ki448=-2;
reg signed [w10-1:0] ka449=65;	reg signed [w10-1:0] kb449=-120;	reg signed [w10-1:0] kc449=44;	reg signed [w10-1:0] kd449=-66;	reg signed [w10-1:0] ke449=2;	reg signed [w10-1:0] kf449=49;	reg signed [w10-1:0] kg449=-150;	reg signed [w10-1:0] kh449=71;	reg signed [w10-1:0] ki449=57;
reg signed [w10-1:0] ka450=36;	reg signed [w10-1:0] kb450=-24;	reg signed [w10-1:0] kc450=-89;	reg signed [w10-1:0] kd450=5;	reg signed [w10-1:0] ke450=79;	reg signed [w10-1:0] kf450=-90;	reg signed [w10-1:0] kg450=0;	reg signed [w10-1:0] kh450=-49;	reg signed [w10-1:0] ki450=-30;
reg signed [w10-1:0] ka451=7;	reg signed [w10-1:0] kb451=61;	reg signed [w10-1:0] kc451=-85;	reg signed [w10-1:0] kd451=46;	reg signed [w10-1:0] ke451=81;	reg signed [w10-1:0] kf451=20;	reg signed [w10-1:0] kg451=35;	reg signed [w10-1:0] kh451=86;	reg signed [w10-1:0] ki451=-101;
reg signed [w10-1:0] ka452=109;	reg signed [w10-1:0] kb452=-33;	reg signed [w10-1:0] kc452=119;	reg signed [w10-1:0] kd452=-36;	reg signed [w10-1:0] ke452=-100;	reg signed [w10-1:0] kf452=84;	reg signed [w10-1:0] kg452=-55;	reg signed [w10-1:0] kh452=-125;	reg signed [w10-1:0] ki452=21;
reg signed [w10-1:0] ka453=-54;	reg signed [w10-1:0] kb453=-53;	reg signed [w10-1:0] kc453=39;	reg signed [w10-1:0] kd453=-103;	reg signed [w10-1:0] ke453=-14;	reg signed [w10-1:0] kf453=-25;	reg signed [w10-1:0] kg453=-82;	reg signed [w10-1:0] kh453=34;	reg signed [w10-1:0] ki453=-23;
reg signed [w10-1:0] ka454=-8;	reg signed [w10-1:0] kb454=73;	reg signed [w10-1:0] kc454=-136;	reg signed [w10-1:0] kd454=125;	reg signed [w10-1:0] ke454=-6;	reg signed [w10-1:0] kf454=96;	reg signed [w10-1:0] kg454=41;	reg signed [w10-1:0] kh454=74;	reg signed [w10-1:0] ki454=83;
reg signed [w10-1:0] ka455=-16;	reg signed [w10-1:0] kb455=118;	reg signed [w10-1:0] kc455=-58;	reg signed [w10-1:0] kd455=54;	reg signed [w10-1:0] ke455=-5;	reg signed [w10-1:0] kf455=-71;	reg signed [w10-1:0] kg455=18;	reg signed [w10-1:0] kh455=27;	reg signed [w10-1:0] ki455=-72;
reg signed [w10-1:0] ka456=-5;	reg signed [w10-1:0] kb456=62;	reg signed [w10-1:0] kc456=20;	reg signed [w10-1:0] kd456=56;	reg signed [w10-1:0] ke456=-21;	reg signed [w10-1:0] kf456=22;	reg signed [w10-1:0] kg456=-92;	reg signed [w10-1:0] kh456=74;	reg signed [w10-1:0] ki456=-117;
reg signed [w10-1:0] ka457=-67;	reg signed [w10-1:0] kb457=6;	reg signed [w10-1:0] kc457=-14;	reg signed [w10-1:0] kd457=-18;	reg signed [w10-1:0] ke457=-116;	reg signed [w10-1:0] kf457=93;	reg signed [w10-1:0] kg457=86;	reg signed [w10-1:0] kh457=89;	reg signed [w10-1:0] ki457=-38;
reg signed [w10-1:0] ka458=75;	reg signed [w10-1:0] kb458=77;	reg signed [w10-1:0] kc458=48;	reg signed [w10-1:0] kd458=-103;	reg signed [w10-1:0] ke458=62;	reg signed [w10-1:0] kf458=25;	reg signed [w10-1:0] kg458=-55;	reg signed [w10-1:0] kh458=106;	reg signed [w10-1:0] ki458=89;
reg signed [w10-1:0] ka459=74;	reg signed [w10-1:0] kb459=59;	reg signed [w10-1:0] kc459=-57;	reg signed [w10-1:0] kd459=112;	reg signed [w10-1:0] ke459=-32;	reg signed [w10-1:0] kf459=-135;	reg signed [w10-1:0] kg459=46;	reg signed [w10-1:0] kh459=-130;	reg signed [w10-1:0] ki459=4;
reg signed [w10-1:0] ka460=120;	reg signed [w10-1:0] kb460=-98;	reg signed [w10-1:0] kc460=-82;	reg signed [w10-1:0] kd460=-33;	reg signed [w10-1:0] ke460=-42;	reg signed [w10-1:0] kf460=27;	reg signed [w10-1:0] kg460=82;	reg signed [w10-1:0] kh460=-59;	reg signed [w10-1:0] ki460=-95;
reg signed [w10-1:0] ka461=95;	reg signed [w10-1:0] kb461=82;	reg signed [w10-1:0] kc461=53;	reg signed [w10-1:0] kd461=-44;	reg signed [w10-1:0] ke461=111;	reg signed [w10-1:0] kf461=74;	reg signed [w10-1:0] kg461=-51;	reg signed [w10-1:0] kh461=126;	reg signed [w10-1:0] ki461=98;
reg signed [w10-1:0] ka462=86;	reg signed [w10-1:0] kb462=-67;	reg signed [w10-1:0] kc462=52;	reg signed [w10-1:0] kd462=-67;	reg signed [w10-1:0] ke462=-26;	reg signed [w10-1:0] kf462=-59;	reg signed [w10-1:0] kg462=6;	reg signed [w10-1:0] kh462=62;	reg signed [w10-1:0] ki462=59;
reg signed [w10-1:0] ka463=94;	reg signed [w10-1:0] kb463=-74;	reg signed [w10-1:0] kc463=46;	reg signed [w10-1:0] kd463=68;	reg signed [w10-1:0] ke463=71;	reg signed [w10-1:0] kf463=-14;	reg signed [w10-1:0] kg463=120;	reg signed [w10-1:0] kh463=107;	reg signed [w10-1:0] ki463=-52;
reg signed [w10-1:0] ka464=-118;	reg signed [w10-1:0] kb464=-29;	reg signed [w10-1:0] kc464=-48;	reg signed [w10-1:0] kd464=-10;	reg signed [w10-1:0] ke464=-16;	reg signed [w10-1:0] kf464=19;	reg signed [w10-1:0] kg464=-68;	reg signed [w10-1:0] kh464=81;	reg signed [w10-1:0] ki464=-49;
reg signed [w10-1:0] ka465=-78;	reg signed [w10-1:0] kb465=-18;	reg signed [w10-1:0] kc465=-28;	reg signed [w10-1:0] kd465=-83;	reg signed [w10-1:0] ke465=72;	reg signed [w10-1:0] kf465=95;	reg signed [w10-1:0] kg465=106;	reg signed [w10-1:0] kh465=66;	reg signed [w10-1:0] ki465=108;
reg signed [w10-1:0] ka466=-3;	reg signed [w10-1:0] kb466=68;	reg signed [w10-1:0] kc466=-76;	reg signed [w10-1:0] kd466=72;	reg signed [w10-1:0] ke466=-116;	reg signed [w10-1:0] kf466=-128;	reg signed [w10-1:0] kg466=0;	reg signed [w10-1:0] kh466=71;	reg signed [w10-1:0] ki466=60;
reg signed [w10-1:0] ka467=-67;	reg signed [w10-1:0] kb467=-77;	reg signed [w10-1:0] kc467=-3;	reg signed [w10-1:0] kd467=50;	reg signed [w10-1:0] ke467=41;	reg signed [w10-1:0] kf467=106;	reg signed [w10-1:0] kg467=88;	reg signed [w10-1:0] kh467=17;	reg signed [w10-1:0] ki467=-93;
reg signed [w10-1:0] ka468=-50;	reg signed [w10-1:0] kb468=-7;	reg signed [w10-1:0] kc468=-22;	reg signed [w10-1:0] kd468=40;	reg signed [w10-1:0] ke468=109;	reg signed [w10-1:0] kf468=76;	reg signed [w10-1:0] kg468=81;	reg signed [w10-1:0] kh468=-81;	reg signed [w10-1:0] ki468=-103;
reg signed [w10-1:0] ka469=-84;	reg signed [w10-1:0] kb469=84;	reg signed [w10-1:0] kc469=-1;	reg signed [w10-1:0] kd469=-88;	reg signed [w10-1:0] ke469=-145;	reg signed [w10-1:0] kf469=126;	reg signed [w10-1:0] kg469=82;	reg signed [w10-1:0] kh469=-56;	reg signed [w10-1:0] ki469=97;
reg signed [w10-1:0] ka470=24;	reg signed [w10-1:0] kb470=-51;	reg signed [w10-1:0] kc470=-30;	reg signed [w10-1:0] kd470=120;	reg signed [w10-1:0] ke470=18;	reg signed [w10-1:0] kf470=61;	reg signed [w10-1:0] kg470=-16;	reg signed [w10-1:0] kh470=-11;	reg signed [w10-1:0] ki470=87;
reg signed [w10-1:0] ka471=25;	reg signed [w10-1:0] kb471=-100;	reg signed [w10-1:0] kc471=-30;	reg signed [w10-1:0] kd471=44;	reg signed [w10-1:0] ke471=-105;	reg signed [w10-1:0] kf471=13;	reg signed [w10-1:0] kg471=-57;	reg signed [w10-1:0] kh471=26;	reg signed [w10-1:0] ki471=65;
reg signed [w10-1:0] ka472=34;	reg signed [w10-1:0] kb472=-61;	reg signed [w10-1:0] kc472=31;	reg signed [w10-1:0] kd472=60;	reg signed [w10-1:0] ke472=-13;	reg signed [w10-1:0] kf472=-124;	reg signed [w10-1:0] kg472=-99;	reg signed [w10-1:0] kh472=64;	reg signed [w10-1:0] ki472=70;
reg signed [w10-1:0] ka473=125;	reg signed [w10-1:0] kb473=164;	reg signed [w10-1:0] kc473=-21;	reg signed [w10-1:0] kd473=32;	reg signed [w10-1:0] ke473=-50;	reg signed [w10-1:0] kf473=-78;	reg signed [w10-1:0] kg473=-82;	reg signed [w10-1:0] kh473=105;	reg signed [w10-1:0] ki473=-106;
reg signed [w10-1:0] ka474=-54;	reg signed [w10-1:0] kb474=-134;	reg signed [w10-1:0] kc474=14;	reg signed [w10-1:0] kd474=-13;	reg signed [w10-1:0] ke474=63;	reg signed [w10-1:0] kf474=-46;	reg signed [w10-1:0] kg474=-8;	reg signed [w10-1:0] kh474=-16;	reg signed [w10-1:0] ki474=54;
reg signed [w10-1:0] ka475=-8;	reg signed [w10-1:0] kb475=117;	reg signed [w10-1:0] kc475=24;	reg signed [w10-1:0] kd475=53;	reg signed [w10-1:0] ke475=-52;	reg signed [w10-1:0] kf475=120;	reg signed [w10-1:0] kg475=-46;	reg signed [w10-1:0] kh475=-66;	reg signed [w10-1:0] ki475=-37;
reg signed [w10-1:0] ka476=-2;	reg signed [w10-1:0] kb476=65;	reg signed [w10-1:0] kc476=-61;	reg signed [w10-1:0] kd476=-140;	reg signed [w10-1:0] ke476=24;	reg signed [w10-1:0] kf476=-55;	reg signed [w10-1:0] kg476=-62;	reg signed [w10-1:0] kh476=20;	reg signed [w10-1:0] ki476=-26;
reg signed [w10-1:0] ka477=61;	reg signed [w10-1:0] kb477=12;	reg signed [w10-1:0] kc477=78;	reg signed [w10-1:0] kd477=-42;	reg signed [w10-1:0] ke477=-76;	reg signed [w10-1:0] kf477=48;	reg signed [w10-1:0] kg477=82;	reg signed [w10-1:0] kh477=-98;	reg signed [w10-1:0] ki477=134;
reg signed [w10-1:0] ka478=-35;	reg signed [w10-1:0] kb478=-82;	reg signed [w10-1:0] kc478=86;	reg signed [w10-1:0] kd478=89;	reg signed [w10-1:0] ke478=-103;	reg signed [w10-1:0] kf478=-63;	reg signed [w10-1:0] kg478=20;	reg signed [w10-1:0] kh478=-89;	reg signed [w10-1:0] ki478=-75;
reg signed [w10-1:0] ka479=-39;	reg signed [w10-1:0] kb479=-92;	reg signed [w10-1:0] kc479=74;	reg signed [w10-1:0] kd479=-68;	reg signed [w10-1:0] ke479=-83;	reg signed [w10-1:0] kf479=-22;	reg signed [w10-1:0] kg479=-10;	reg signed [w10-1:0] kh479=50;	reg signed [w10-1:0] ki479=-39;
reg signed [w10-1:0] ka480=89;	reg signed [w10-1:0] kb480=-70;	reg signed [w10-1:0] kc480=-47;	reg signed [w10-1:0] kd480=22;	reg signed [w10-1:0] ke480=-92;	reg signed [w10-1:0] kf480=29;	reg signed [w10-1:0] kg480=-10;	reg signed [w10-1:0] kh480=148;	reg signed [w10-1:0] ki480=24;
reg signed [w10-1:0] ka481=88;	reg signed [w10-1:0] kb481=-73;	reg signed [w10-1:0] kc481=-5;	reg signed [w10-1:0] kd481=-95;	reg signed [w10-1:0] ke481=-106;	reg signed [w10-1:0] kf481=113;	reg signed [w10-1:0] kg481=-83;	reg signed [w10-1:0] kh481=41;	reg signed [w10-1:0] ki481=-32;
reg signed [w10-1:0] ka482=100;	reg signed [w10-1:0] kb482=-11;	reg signed [w10-1:0] kc482=-8;	reg signed [w10-1:0] kd482=27;	reg signed [w10-1:0] ke482=-29;	reg signed [w10-1:0] kf482=-8;	reg signed [w10-1:0] kg482=117;	reg signed [w10-1:0] kh482=-11;	reg signed [w10-1:0] ki482=136;
reg signed [w10-1:0] ka483=75;	reg signed [w10-1:0] kb483=79;	reg signed [w10-1:0] kc483=-102;	reg signed [w10-1:0] kd483=-41;	reg signed [w10-1:0] ke483=-57;	reg signed [w10-1:0] kf483=64;	reg signed [w10-1:0] kg483=68;	reg signed [w10-1:0] kh483=-77;	reg signed [w10-1:0] ki483=23;
reg signed [w10-1:0] ka484=27;	reg signed [w10-1:0] kb484=-32;	reg signed [w10-1:0] kc484=-64;	reg signed [w10-1:0] kd484=77;	reg signed [w10-1:0] ke484=54;	reg signed [w10-1:0] kf484=-64;	reg signed [w10-1:0] kg484=-49;	reg signed [w10-1:0] kh484=-20;	reg signed [w10-1:0] ki484=-2;
reg signed [w10-1:0] ka485=95;	reg signed [w10-1:0] kb485=27;	reg signed [w10-1:0] kc485=-35;	reg signed [w10-1:0] kd485=-102;	reg signed [w10-1:0] ke485=98;	reg signed [w10-1:0] kf485=-117;	reg signed [w10-1:0] kg485=-76;	reg signed [w10-1:0] kh485=-43;	reg signed [w10-1:0] ki485=-121;
reg signed [w10-1:0] ka486=5;	reg signed [w10-1:0] kb486=-39;	reg signed [w10-1:0] kc486=54;	reg signed [w10-1:0] kd486=82;	reg signed [w10-1:0] ke486=-89;	reg signed [w10-1:0] kf486=-116;	reg signed [w10-1:0] kg486=-20;	reg signed [w10-1:0] kh486=-7;	reg signed [w10-1:0] ki486=-59;
reg signed [w10-1:0] ka487=75;	reg signed [w10-1:0] kb487=94;	reg signed [w10-1:0] kc487=96;	reg signed [w10-1:0] kd487=-108;	reg signed [w10-1:0] ke487=101;	reg signed [w10-1:0] kf487=25;	reg signed [w10-1:0] kg487=26;	reg signed [w10-1:0] kh487=18;	reg signed [w10-1:0] ki487=103;
reg signed [w10-1:0] ka488=-43;	reg signed [w10-1:0] kb488=72;	reg signed [w10-1:0] kc488=-96;	reg signed [w10-1:0] kd488=-76;	reg signed [w10-1:0] ke488=7;	reg signed [w10-1:0] kf488=-7;	reg signed [w10-1:0] kg488=60;	reg signed [w10-1:0] kh488=-3;	reg signed [w10-1:0] ki488=1;
reg signed [w10-1:0] ka489=-28;	reg signed [w10-1:0] kb489=19;	reg signed [w10-1:0] kc489=155;	reg signed [w10-1:0] kd489=143;	reg signed [w10-1:0] ke489=68;	reg signed [w10-1:0] kf489=112;	reg signed [w10-1:0] kg489=71;	reg signed [w10-1:0] kh489=56;	reg signed [w10-1:0] ki489=80;
reg signed [w10-1:0] ka490=72;	reg signed [w10-1:0] kb490=86;	reg signed [w10-1:0] kc490=15;	reg signed [w10-1:0] kd490=-146;	reg signed [w10-1:0] ke490=-14;	reg signed [w10-1:0] kf490=-89;	reg signed [w10-1:0] kg490=34;	reg signed [w10-1:0] kh490=-104;	reg signed [w10-1:0] ki490=-35;
reg signed [w10-1:0] ka491=-100;	reg signed [w10-1:0] kb491=-44;	reg signed [w10-1:0] kc491=-84;	reg signed [w10-1:0] kd491=-91;	reg signed [w10-1:0] ke491=5;	reg signed [w10-1:0] kf491=95;	reg signed [w10-1:0] kg491=111;	reg signed [w10-1:0] kh491=14;	reg signed [w10-1:0] ki491=-16;
reg signed [w10-1:0] ka492=100;	reg signed [w10-1:0] kb492=-22;	reg signed [w10-1:0] kc492=-55;	reg signed [w10-1:0] kd492=-103;	reg signed [w10-1:0] ke492=-62;	reg signed [w10-1:0] kf492=-68;	reg signed [w10-1:0] kg492=127;	reg signed [w10-1:0] kh492=-30;	reg signed [w10-1:0] ki492=107;
reg signed [w10-1:0] ka493=88;	reg signed [w10-1:0] kb493=-123;	reg signed [w10-1:0] kc493=62;	reg signed [w10-1:0] kd493=86;	reg signed [w10-1:0] ke493=92;	reg signed [w10-1:0] kf493=-45;	reg signed [w10-1:0] kg493=-88;	reg signed [w10-1:0] kh493=3;	reg signed [w10-1:0] ki493=-84;
reg signed [w10-1:0] ka494=-26;	reg signed [w10-1:0] kb494=-95;	reg signed [w10-1:0] kc494=153;	reg signed [w10-1:0] kd494=-27;	reg signed [w10-1:0] ke494=-74;	reg signed [w10-1:0] kf494=46;	reg signed [w10-1:0] kg494=99;	reg signed [w10-1:0] kh494=-63;	reg signed [w10-1:0] ki494=-116;
reg signed [w10-1:0] ka495=57;	reg signed [w10-1:0] kb495=114;	reg signed [w10-1:0] kc495=42;	reg signed [w10-1:0] kd495=-27;	reg signed [w10-1:0] ke495=43;	reg signed [w10-1:0] kf495=-77;	reg signed [w10-1:0] kg495=33;	reg signed [w10-1:0] kh495=-50;	reg signed [w10-1:0] ki495=-93;
reg signed [w10-1:0] ka496=-75;	reg signed [w10-1:0] kb496=-23;	reg signed [w10-1:0] kc496=105;	reg signed [w10-1:0] kd496=-34;	reg signed [w10-1:0] ke496=-99;	reg signed [w10-1:0] kf496=-59;	reg signed [w10-1:0] kg496=68;	reg signed [w10-1:0] kh496=-74;	reg signed [w10-1:0] ki496=-74;
reg signed [w10-1:0] ka497=89;	reg signed [w10-1:0] kb497=-84;	reg signed [w10-1:0] kc497=16;	reg signed [w10-1:0] kd497=-81;	reg signed [w10-1:0] ke497=-37;	reg signed [w10-1:0] kf497=40;	reg signed [w10-1:0] kg497=63;	reg signed [w10-1:0] kh497=69;	reg signed [w10-1:0] ki497=69;
reg signed [w10-1:0] ka498=-34;	reg signed [w10-1:0] kb498=50;	reg signed [w10-1:0] kc498=-48;	reg signed [w10-1:0] kd498=-55;	reg signed [w10-1:0] ke498=-28;	reg signed [w10-1:0] kf498=67;	reg signed [w10-1:0] kg498=-27;	reg signed [w10-1:0] kh498=133;	reg signed [w10-1:0] ki498=68;
reg signed [w10-1:0] ka499=-24;	reg signed [w10-1:0] kb499=124;	reg signed [w10-1:0] kc499=-7;	reg signed [w10-1:0] kd499=63;	reg signed [w10-1:0] ke499=56;	reg signed [w10-1:0] kf499=-53;	reg signed [w10-1:0] kg499=13;	reg signed [w10-1:0] kh499=114;	reg signed [w10-1:0] ki499=42;
reg signed [w10-1:0] ka500=42;	reg signed [w10-1:0] kb500=2;	reg signed [w10-1:0] kc500=-64;	reg signed [w10-1:0] kd500=12;	reg signed [w10-1:0] ke500=-65;	reg signed [w10-1:0] kf500=32;	reg signed [w10-1:0] kg500=-24;	reg signed [w10-1:0] kh500=93;	reg signed [w10-1:0] ki500=-35;
reg signed [w10-1:0] ka501=77;	reg signed [w10-1:0] kb501=119;	reg signed [w10-1:0] kc501=119;	reg signed [w10-1:0] kd501=83;	reg signed [w10-1:0] ke501=47;	reg signed [w10-1:0] kf501=120;	reg signed [w10-1:0] kg501=35;	reg signed [w10-1:0] kh501=20;	reg signed [w10-1:0] ki501=81;
reg signed [w10-1:0] ka502=9;	reg signed [w10-1:0] kb502=-15;	reg signed [w10-1:0] kc502=112;	reg signed [w10-1:0] kd502=23;	reg signed [w10-1:0] ke502=102;	reg signed [w10-1:0] kf502=-81;	reg signed [w10-1:0] kg502=-98;	reg signed [w10-1:0] kh502=-62;	reg signed [w10-1:0] ki502=-35;
reg signed [w10-1:0] ka503=-87;	reg signed [w10-1:0] kb503=-99;	reg signed [w10-1:0] kc503=25;	reg signed [w10-1:0] kd503=24;	reg signed [w10-1:0] ke503=71;	reg signed [w10-1:0] kf503=-11;	reg signed [w10-1:0] kg503=82;	reg signed [w10-1:0] kh503=5;	reg signed [w10-1:0] ki503=125;
reg signed [w10-1:0] ka504=127;	reg signed [w10-1:0] kb504=-5;	reg signed [w10-1:0] kc504=-24;	reg signed [w10-1:0] kd504=11;	reg signed [w10-1:0] ke504=41;	reg signed [w10-1:0] kf504=-20;	reg signed [w10-1:0] kg504=-74;	reg signed [w10-1:0] kh504=21;	reg signed [w10-1:0] ki504=-131;
reg signed [w10-1:0] ka505=-39;	reg signed [w10-1:0] kb505=-9;	reg signed [w10-1:0] kc505=103;	reg signed [w10-1:0] kd505=-97;	reg signed [w10-1:0] ke505=-114;	reg signed [w10-1:0] kf505=-105;	reg signed [w10-1:0] kg505=-77;	reg signed [w10-1:0] kh505=-138;	reg signed [w10-1:0] ki505=-61;
reg signed [w10-1:0] ka506=93;	reg signed [w10-1:0] kb506=15;	reg signed [w10-1:0] kc506=-105;	reg signed [w10-1:0] kd506=39;	reg signed [w10-1:0] ke506=-4;	reg signed [w10-1:0] kf506=43;	reg signed [w10-1:0] kg506=122;	reg signed [w10-1:0] kh506=-23;	reg signed [w10-1:0] ki506=48;
reg signed [w10-1:0] ka507=11;	reg signed [w10-1:0] kb507=-176;	reg signed [w10-1:0] kc507=67;	reg signed [w10-1:0] kd507=45;	reg signed [w10-1:0] ke507=-21;	reg signed [w10-1:0] kf507=-19;	reg signed [w10-1:0] kg507=-37;	reg signed [w10-1:0] kh507=38;	reg signed [w10-1:0] ki507=-93;
reg signed [w10-1:0] ka508=-59;	reg signed [w10-1:0] kb508=-63;	reg signed [w10-1:0] kc508=6;	reg signed [w10-1:0] kd508=-99;	reg signed [w10-1:0] ke508=-45;	reg signed [w10-1:0] kf508=87;	reg signed [w10-1:0] kg508=-27;	reg signed [w10-1:0] kh508=-85;	reg signed [w10-1:0] ki508=-82;
reg signed [w10-1:0] ka509=-64;	reg signed [w10-1:0] kb509=-41;	reg signed [w10-1:0] kc509=99;	reg signed [w10-1:0] kd509=-72;	reg signed [w10-1:0] ke509=-56;	reg signed [w10-1:0] kf509=70;	reg signed [w10-1:0] kg509=114;	reg signed [w10-1:0] kh509=87;	reg signed [w10-1:0] ki509=-24;
reg signed [w10-1:0] ka510=-22;	reg signed [w10-1:0] kb510=100;	reg signed [w10-1:0] kc510=-33;	reg signed [w10-1:0] kd510=85;	reg signed [w10-1:0] ke510=61;	reg signed [w10-1:0] kf510=66;	reg signed [w10-1:0] kg510=-40;	reg signed [w10-1:0] kh510=46;	reg signed [w10-1:0] ki510=143;
reg signed [w10-1:0] ka511=-84;	reg signed [w10-1:0] kb511=-11;	reg signed [w10-1:0] kc511=53;	reg signed [w10-1:0] kd511=108;	reg signed [w10-1:0] ke511=43;	reg signed [w10-1:0] kf511=88;	reg signed [w10-1:0] kg511=57;	reg signed [w10-1:0] kh511=96;	reg signed [w10-1:0] ki511=-103;
reg signed [w10-1:0] ka512=-58;	reg signed [w10-1:0] kb512=76;	reg signed [w10-1:0] kc512=35;	reg signed [w10-1:0] kd512=-39;	reg signed [w10-1:0] ke512=114;	reg signed [w10-1:0] kf512=107;	reg signed [w10-1:0] kg512=28;	reg signed [w10-1:0] kh512=33;	reg signed [w10-1:0] ki512=17;
reg signed [w10-1:0] ka513=82;	reg signed [w10-1:0] kb513=-64;	reg signed [w10-1:0] kc513=-8;	reg signed [w10-1:0] kd513=-71;	reg signed [w10-1:0] ke513=94;	reg signed [w10-1:0] kf513=-45;	reg signed [w10-1:0] kg513=-20;	reg signed [w10-1:0] kh513=-32;	reg signed [w10-1:0] ki513=-99;
reg signed [w10-1:0] ka514=128;	reg signed [w10-1:0] kb514=-40;	reg signed [w10-1:0] kc514=-125;	reg signed [w10-1:0] kd514=-103;	reg signed [w10-1:0] ke514=-132;	reg signed [w10-1:0] kf514=-140;	reg signed [w10-1:0] kg514=100;	reg signed [w10-1:0] kh514=12;	reg signed [w10-1:0] ki514=39;
reg signed [w10-1:0] ka515=-138;	reg signed [w10-1:0] kb515=-59;	reg signed [w10-1:0] kc515=7;	reg signed [w10-1:0] kd515=-114;	reg signed [w10-1:0] ke515=8;	reg signed [w10-1:0] kf515=-19;	reg signed [w10-1:0] kg515=-66;	reg signed [w10-1:0] kh515=-3;	reg signed [w10-1:0] ki515=-95;
reg signed [w10-1:0] ka516=-2;	reg signed [w10-1:0] kb516=-18;	reg signed [w10-1:0] kc516=-61;	reg signed [w10-1:0] kd516=-3;	reg signed [w10-1:0] ke516=16;	reg signed [w10-1:0] kf516=-11;	reg signed [w10-1:0] kg516=-103;	reg signed [w10-1:0] kh516=-108;	reg signed [w10-1:0] ki516=-63;
reg signed [w10-1:0] ka517=-32;	reg signed [w10-1:0] kb517=11;	reg signed [w10-1:0] kc517=-24;	reg signed [w10-1:0] kd517=-69;	reg signed [w10-1:0] ke517=-18;	reg signed [w10-1:0] kf517=110;	reg signed [w10-1:0] kg517=-38;	reg signed [w10-1:0] kh517=84;	reg signed [w10-1:0] ki517=22;
reg signed [w10-1:0] ka518=13;	reg signed [w10-1:0] kb518=-1;	reg signed [w10-1:0] kc518=53;	reg signed [w10-1:0] kd518=57;	reg signed [w10-1:0] ke518=29;	reg signed [w10-1:0] kf518=-124;	reg signed [w10-1:0] kg518=-11;	reg signed [w10-1:0] kh518=14;	reg signed [w10-1:0] ki518=-49;
reg signed [w10-1:0] ka519=-56;	reg signed [w10-1:0] kb519=-62;	reg signed [w10-1:0] kc519=-123;	reg signed [w10-1:0] kd519=-32;	reg signed [w10-1:0] ke519=-121;	reg signed [w10-1:0] kf519=3;	reg signed [w10-1:0] kg519=-90;	reg signed [w10-1:0] kh519=-172;	reg signed [w10-1:0] ki519=-76;
reg signed [w10-1:0] ka520=82;	reg signed [w10-1:0] kb520=31;	reg signed [w10-1:0] kc520=54;	reg signed [w10-1:0] kd520=-24;	reg signed [w10-1:0] ke520=95;	reg signed [w10-1:0] kf520=19;	reg signed [w10-1:0] kg520=82;	reg signed [w10-1:0] kh520=-56;	reg signed [w10-1:0] ki520=7;
reg signed [w10-1:0] ka521=-7;	reg signed [w10-1:0] kb521=35;	reg signed [w10-1:0] kc521=38;	reg signed [w10-1:0] kd521=85;	reg signed [w10-1:0] ke521=42;	reg signed [w10-1:0] kf521=56;	reg signed [w10-1:0] kg521=58;	reg signed [w10-1:0] kh521=-110;	reg signed [w10-1:0] ki521=73;
reg signed [w10-1:0] ka522=-8;	reg signed [w10-1:0] kb522=-117;	reg signed [w10-1:0] kc522=70;	reg signed [w10-1:0] kd522=97;	reg signed [w10-1:0] ke522=-84;	reg signed [w10-1:0] kf522=-70;	reg signed [w10-1:0] kg522=-51;	reg signed [w10-1:0] kh522=93;	reg signed [w10-1:0] ki522=-69;
reg signed [w10-1:0] ka523=45;	reg signed [w10-1:0] kb523=23;	reg signed [w10-1:0] kc523=-33;	reg signed [w10-1:0] kd523=-20;	reg signed [w10-1:0] ke523=-24;	reg signed [w10-1:0] kf523=-14;	reg signed [w10-1:0] kg523=132;	reg signed [w10-1:0] kh523=-59;	reg signed [w10-1:0] ki523=-52;
reg signed [w10-1:0] ka524=138;	reg signed [w10-1:0] kb524=97;	reg signed [w10-1:0] kc524=-50;	reg signed [w10-1:0] kd524=-48;	reg signed [w10-1:0] ke524=-84;	reg signed [w10-1:0] kf524=-116;	reg signed [w10-1:0] kg524=39;	reg signed [w10-1:0] kh524=27;	reg signed [w10-1:0] ki524=-31;
reg signed [w10-1:0] ka525=-134;	reg signed [w10-1:0] kb525=-81;	reg signed [w10-1:0] kc525=39;	reg signed [w10-1:0] kd525=-49;	reg signed [w10-1:0] ke525=-118;	reg signed [w10-1:0] kf525=112;	reg signed [w10-1:0] kg525=10;	reg signed [w10-1:0] kh525=86;	reg signed [w10-1:0] ki525=103;
reg signed [w10-1:0] ka526=3;	reg signed [w10-1:0] kb526=-49;	reg signed [w10-1:0] kc526=-106;	reg signed [w10-1:0] kd526=120;	reg signed [w10-1:0] ke526=63;	reg signed [w10-1:0] kf526=-131;	reg signed [w10-1:0] kg526=83;	reg signed [w10-1:0] kh526=-85;	reg signed [w10-1:0] ki526=-62;
reg signed [w10-1:0] ka527=-53;	reg signed [w10-1:0] kb527=94;	reg signed [w10-1:0] kc527=24;	reg signed [w10-1:0] kd527=-107;	reg signed [w10-1:0] ke527=-7;	reg signed [w10-1:0] kf527=-77;	reg signed [w10-1:0] kg527=55;	reg signed [w10-1:0] kh527=99;	reg signed [w10-1:0] ki527=79;
reg signed [w10-1:0] ka528=92;	reg signed [w10-1:0] kb528=30;	reg signed [w10-1:0] kc528=-76;	reg signed [w10-1:0] kd528=-119;	reg signed [w10-1:0] ke528=146;	reg signed [w10-1:0] kf528=-97;	reg signed [w10-1:0] kg528=-52;	reg signed [w10-1:0] kh528=133;	reg signed [w10-1:0] ki528=-114;
reg signed [w10-1:0] ka529=34;	reg signed [w10-1:0] kb529=-31;	reg signed [w10-1:0] kc529=21;	reg signed [w10-1:0] kd529=-29;	reg signed [w10-1:0] ke529=-73;	reg signed [w10-1:0] kf529=21;	reg signed [w10-1:0] kg529=-53;	reg signed [w10-1:0] kh529=110;	reg signed [w10-1:0] ki529=78;
reg signed [w10-1:0] ka530=-47;	reg signed [w10-1:0] kb530=-58;	reg signed [w10-1:0] kc530=-53;	reg signed [w10-1:0] kd530=20;	reg signed [w10-1:0] ke530=20;	reg signed [w10-1:0] kf530=5;	reg signed [w10-1:0] kg530=108;	reg signed [w10-1:0] kh530=117;	reg signed [w10-1:0] ki530=-17;
reg signed [w10-1:0] ka531=98;	reg signed [w10-1:0] kb531=20;	reg signed [w10-1:0] kc531=-13;	reg signed [w10-1:0] kd531=-115;	reg signed [w10-1:0] ke531=2;	reg signed [w10-1:0] kf531=-38;	reg signed [w10-1:0] kg531=44;	reg signed [w10-1:0] kh531=64;	reg signed [w10-1:0] ki531=20;
reg signed [w10-1:0] ka532=11;	reg signed [w10-1:0] kb532=-54;	reg signed [w10-1:0] kc532=-11;	reg signed [w10-1:0] kd532=-56;	reg signed [w10-1:0] ke532=109;	reg signed [w10-1:0] kf532=-65;	reg signed [w10-1:0] kg532=-152;	reg signed [w10-1:0] kh532=109;	reg signed [w10-1:0] ki532=-7;
reg signed [w10-1:0] ka533=121;	reg signed [w10-1:0] kb533=78;	reg signed [w10-1:0] kc533=-25;	reg signed [w10-1:0] kd533=1;	reg signed [w10-1:0] ke533=-63;	reg signed [w10-1:0] kf533=-103;	reg signed [w10-1:0] kg533=74;	reg signed [w10-1:0] kh533=-75;	reg signed [w10-1:0] ki533=49;
reg signed [w10-1:0] ka534=-49;	reg signed [w10-1:0] kb534=48;	reg signed [w10-1:0] kc534=-41;	reg signed [w10-1:0] kd534=-7;	reg signed [w10-1:0] ke534=-64;	reg signed [w10-1:0] kf534=4;	reg signed [w10-1:0] kg534=-72;	reg signed [w10-1:0] kh534=52;	reg signed [w10-1:0] ki534=-66;
reg signed [w10-1:0] ka535=81;	reg signed [w10-1:0] kb535=-72;	reg signed [w10-1:0] kc535=-49;	reg signed [w10-1:0] kd535=-89;	reg signed [w10-1:0] ke535=-23;	reg signed [w10-1:0] kf535=59;	reg signed [w10-1:0] kg535=-69;	reg signed [w10-1:0] kh535=-32;	reg signed [w10-1:0] ki535=101;
reg signed [w10-1:0] ka536=-29;	reg signed [w10-1:0] kb536=177;	reg signed [w10-1:0] kc536=91;	reg signed [w10-1:0] kd536=113;	reg signed [w10-1:0] ke536=-39;	reg signed [w10-1:0] kf536=44;	reg signed [w10-1:0] kg536=108;	reg signed [w10-1:0] kh536=-55;	reg signed [w10-1:0] ki536=150;
reg signed [w10-1:0] ka537=52;	reg signed [w10-1:0] kb537=2;	reg signed [w10-1:0] kc537=-6;	reg signed [w10-1:0] kd537=36;	reg signed [w10-1:0] ke537=51;	reg signed [w10-1:0] kf537=5;	reg signed [w10-1:0] kg537=-8;	reg signed [w10-1:0] kh537=65;	reg signed [w10-1:0] ki537=-125;
reg signed [w10-1:0] ka538=-55;	reg signed [w10-1:0] kb538=-126;	reg signed [w10-1:0] kc538=46;	reg signed [w10-1:0] kd538=122;	reg signed [w10-1:0] ke538=-55;	reg signed [w10-1:0] kf538=36;	reg signed [w10-1:0] kg538=30;	reg signed [w10-1:0] kh538=-125;	reg signed [w10-1:0] ki538=-14;
reg signed [w10-1:0] ka539=70;	reg signed [w10-1:0] kb539=25;	reg signed [w10-1:0] kc539=-12;	reg signed [w10-1:0] kd539=-26;	reg signed [w10-1:0] ke539=68;	reg signed [w10-1:0] kf539=37;	reg signed [w10-1:0] kg539=-45;	reg signed [w10-1:0] kh539=30;	reg signed [w10-1:0] ki539=1;
reg signed [w10-1:0] ka540=-119;	reg signed [w10-1:0] kb540=-69;	reg signed [w10-1:0] kc540=-118;	reg signed [w10-1:0] kd540=97;	reg signed [w10-1:0] ke540=-79;	reg signed [w10-1:0] kf540=100;	reg signed [w10-1:0] kg540=157;	reg signed [w10-1:0] kh540=-66;	reg signed [w10-1:0] ki540=73;
reg signed [w10-1:0] ka541=11;	reg signed [w10-1:0] kb541=116;	reg signed [w10-1:0] kc541=-24;	reg signed [w10-1:0] kd541=-55;	reg signed [w10-1:0] ke541=14;	reg signed [w10-1:0] kf541=58;	reg signed [w10-1:0] kg541=10;	reg signed [w10-1:0] kh541=-103;	reg signed [w10-1:0] ki541=-17;
reg signed [w10-1:0] ka542=115;	reg signed [w10-1:0] kb542=18;	reg signed [w10-1:0] kc542=-95;	reg signed [w10-1:0] kd542=45;	reg signed [w10-1:0] ke542=-1;	reg signed [w10-1:0] kf542=-61;	reg signed [w10-1:0] kg542=77;	reg signed [w10-1:0] kh542=109;	reg signed [w10-1:0] ki542=145;
reg signed [w10-1:0] ka543=48;	reg signed [w10-1:0] kb543=118;	reg signed [w10-1:0] kc543=67;	reg signed [w10-1:0] kd543=-69;	reg signed [w10-1:0] ke543=77;	reg signed [w10-1:0] kf543=-57;	reg signed [w10-1:0] kg543=62;	reg signed [w10-1:0] kh543=27;	reg signed [w10-1:0] ki543=119;
reg signed [w10-1:0] ka544=38;	reg signed [w10-1:0] kb544=-110;	reg signed [w10-1:0] kc544=-65;	reg signed [w10-1:0] kd544=-14;	reg signed [w10-1:0] ke544=-132;	reg signed [w10-1:0] kf544=45;	reg signed [w10-1:0] kg544=146;	reg signed [w10-1:0] kh544=-127;	reg signed [w10-1:0] ki544=-17;
reg signed [w10-1:0] ka545=58;	reg signed [w10-1:0] kb545=48;	reg signed [w10-1:0] kc545=-62;	reg signed [w10-1:0] kd545=22;	reg signed [w10-1:0] ke545=-7;	reg signed [w10-1:0] kf545=-87;	reg signed [w10-1:0] kg545=-121;	reg signed [w10-1:0] kh545=-44;	reg signed [w10-1:0] ki545=-20;
reg signed [w10-1:0] ka546=9;	reg signed [w10-1:0] kb546=50;	reg signed [w10-1:0] kc546=94;	reg signed [w10-1:0] kd546=131;	reg signed [w10-1:0] ke546=-46;	reg signed [w10-1:0] kf546=-52;	reg signed [w10-1:0] kg546=-58;	reg signed [w10-1:0] kh546=123;	reg signed [w10-1:0] ki546=119;
reg signed [w10-1:0] ka547=-76;	reg signed [w10-1:0] kb547=14;	reg signed [w10-1:0] kc547=116;	reg signed [w10-1:0] kd547=103;	reg signed [w10-1:0] ke547=-10;	reg signed [w10-1:0] kf547=75;	reg signed [w10-1:0] kg547=126;	reg signed [w10-1:0] kh547=-75;	reg signed [w10-1:0] ki547=98;
reg signed [w10-1:0] ka548=-44;	reg signed [w10-1:0] kb548=-90;	reg signed [w10-1:0] kc548=-16;	reg signed [w10-1:0] kd548=-120;	reg signed [w10-1:0] ke548=-6;	reg signed [w10-1:0] kf548=-17;	reg signed [w10-1:0] kg548=-143;	reg signed [w10-1:0] kh548=-23;	reg signed [w10-1:0] ki548=75;
reg signed [w10-1:0] ka549=-90;	reg signed [w10-1:0] kb549=101;	reg signed [w10-1:0] kc549=-9;	reg signed [w10-1:0] kd549=7;	reg signed [w10-1:0] ke549=38;	reg signed [w10-1:0] kf549=-15;	reg signed [w10-1:0] kg549=-100;	reg signed [w10-1:0] kh549=12;	reg signed [w10-1:0] ki549=3;
reg signed [w10-1:0] ka550=-26;	reg signed [w10-1:0] kb550=7;	reg signed [w10-1:0] kc550=33;	reg signed [w10-1:0] kd550=151;	reg signed [w10-1:0] ke550=-42;	reg signed [w10-1:0] kf550=-37;	reg signed [w10-1:0] kg550=54;	reg signed [w10-1:0] kh550=-108;	reg signed [w10-1:0] ki550=-5;
reg signed [w10-1:0] ka551=-41;	reg signed [w10-1:0] kb551=146;	reg signed [w10-1:0] kc551=61;	reg signed [w10-1:0] kd551=86;	reg signed [w10-1:0] ke551=-67;	reg signed [w10-1:0] kf551=75;	reg signed [w10-1:0] kg551=-12;	reg signed [w10-1:0] kh551=50;	reg signed [w10-1:0] ki551=-11;
reg signed [w10-1:0] ka552=-85;	reg signed [w10-1:0] kb552=77;	reg signed [w10-1:0] kc552=22;	reg signed [w10-1:0] kd552=-33;	reg signed [w10-1:0] ke552=-83;	reg signed [w10-1:0] kf552=-153;	reg signed [w10-1:0] kg552=87;	reg signed [w10-1:0] kh552=3;	reg signed [w10-1:0] ki552=-15;
reg signed [w10-1:0] ka553=-73;	reg signed [w10-1:0] kb553=7;	reg signed [w10-1:0] kc553=-37;	reg signed [w10-1:0] kd553=69;	reg signed [w10-1:0] ke553=80;	reg signed [w10-1:0] kf553=49;	reg signed [w10-1:0] kg553=141;	reg signed [w10-1:0] kh553=9;	reg signed [w10-1:0] ki553=41;
reg signed [w10-1:0] ka554=5;	reg signed [w10-1:0] kb554=43;	reg signed [w10-1:0] kc554=69;	reg signed [w10-1:0] kd554=-26;	reg signed [w10-1:0] ke554=-74;	reg signed [w10-1:0] kf554=27;	reg signed [w10-1:0] kg554=-99;	reg signed [w10-1:0] kh554=40;	reg signed [w10-1:0] ki554=42;
reg signed [w10-1:0] ka555=44;	reg signed [w10-1:0] kb555=-87;	reg signed [w10-1:0] kc555=-89;	reg signed [w10-1:0] kd555=103;	reg signed [w10-1:0] ke555=132;	reg signed [w10-1:0] kf555=-84;	reg signed [w10-1:0] kg555=-7;	reg signed [w10-1:0] kh555=-126;	reg signed [w10-1:0] ki555=31;
reg signed [w10-1:0] ka556=-128;	reg signed [w10-1:0] kb556=-72;	reg signed [w10-1:0] kc556=111;	reg signed [w10-1:0] kd556=-14;	reg signed [w10-1:0] ke556=55;	reg signed [w10-1:0] kf556=88;	reg signed [w10-1:0] kg556=-13;	reg signed [w10-1:0] kh556=63;	reg signed [w10-1:0] ki556=91;
reg signed [w10-1:0] ka557=-78;	reg signed [w10-1:0] kb557=-2;	reg signed [w10-1:0] kc557=115;	reg signed [w10-1:0] kd557=-127;	reg signed [w10-1:0] ke557=-24;	reg signed [w10-1:0] kf557=11;	reg signed [w10-1:0] kg557=80;	reg signed [w10-1:0] kh557=-53;	reg signed [w10-1:0] ki557=50;
reg signed [w10-1:0] ka558=30;	reg signed [w10-1:0] kb558=-48;	reg signed [w10-1:0] kc558=-15;	reg signed [w10-1:0] kd558=-96;	reg signed [w10-1:0] ke558=75;	reg signed [w10-1:0] kf558=-32;	reg signed [w10-1:0] kg558=25;	reg signed [w10-1:0] kh558=82;	reg signed [w10-1:0] ki558=141;
reg signed [w10-1:0] ka559=-29;	reg signed [w10-1:0] kb559=-44;	reg signed [w10-1:0] kc559=90;	reg signed [w10-1:0] kd559=-35;	reg signed [w10-1:0] ke559=-2;	reg signed [w10-1:0] kf559=45;	reg signed [w10-1:0] kg559=-87;	reg signed [w10-1:0] kh559=45;	reg signed [w10-1:0] ki559=-73;
reg signed [w10-1:0] ka560=118;	reg signed [w10-1:0] kb560=-37;	reg signed [w10-1:0] kc560=67;	reg signed [w10-1:0] kd560=59;	reg signed [w10-1:0] ke560=-120;	reg signed [w10-1:0] kf560=-38;	reg signed [w10-1:0] kg560=-37;	reg signed [w10-1:0] kh560=-54;	reg signed [w10-1:0] ki560=-31;
reg signed [w10-1:0] ka561=105;	reg signed [w10-1:0] kb561=-82;	reg signed [w10-1:0] kc561=-50;	reg signed [w10-1:0] kd561=-6;	reg signed [w10-1:0] ke561=58;	reg signed [w10-1:0] kf561=-94;	reg signed [w10-1:0] kg561=-5;	reg signed [w10-1:0] kh561=-6;	reg signed [w10-1:0] ki561=-72;
reg signed [w10-1:0] ka562=-105;	reg signed [w10-1:0] kb562=-84;	reg signed [w10-1:0] kc562=-37;	reg signed [w10-1:0] kd562=-52;	reg signed [w10-1:0] ke562=49;	reg signed [w10-1:0] kf562=-45;	reg signed [w10-1:0] kg562=-121;	reg signed [w10-1:0] kh562=98;	reg signed [w10-1:0] ki562=-35;
reg signed [w10-1:0] ka563=53;	reg signed [w10-1:0] kb563=-46;	reg signed [w10-1:0] kc563=87;	reg signed [w10-1:0] kd563=-60;	reg signed [w10-1:0] ke563=118;	reg signed [w10-1:0] kf563=146;	reg signed [w10-1:0] kg563=34;	reg signed [w10-1:0] kh563=23;	reg signed [w10-1:0] ki563=106;
reg signed [w10-1:0] ka564=-13;	reg signed [w10-1:0] kb564=16;	reg signed [w10-1:0] kc564=92;	reg signed [w10-1:0] kd564=-71;	reg signed [w10-1:0] ke564=3;	reg signed [w10-1:0] kf564=83;	reg signed [w10-1:0] kg564=-85;	reg signed [w10-1:0] kh564=74;	reg signed [w10-1:0] ki564=-129;
reg signed [w10-1:0] ka565=2;	reg signed [w10-1:0] kb565=7;	reg signed [w10-1:0] kc565=-99;	reg signed [w10-1:0] kd565=115;	reg signed [w10-1:0] ke565=-57;	reg signed [w10-1:0] kf565=82;	reg signed [w10-1:0] kg565=26;	reg signed [w10-1:0] kh565=-48;	reg signed [w10-1:0] ki565=5;
reg signed [w10-1:0] ka566=119;	reg signed [w10-1:0] kb566=61;	reg signed [w10-1:0] kc566=25;	reg signed [w10-1:0] kd566=1;	reg signed [w10-1:0] ke566=-125;	reg signed [w10-1:0] kf566=-66;	reg signed [w10-1:0] kg566=94;	reg signed [w10-1:0] kh566=131;	reg signed [w10-1:0] ki566=134;
reg signed [w10-1:0] ka567=121;	reg signed [w10-1:0] kb567=-35;	reg signed [w10-1:0] kc567=104;	reg signed [w10-1:0] kd567=89;	reg signed [w10-1:0] ke567=138;	reg signed [w10-1:0] kf567=79;	reg signed [w10-1:0] kg567=11;	reg signed [w10-1:0] kh567=54;	reg signed [w10-1:0] ki567=-45;
reg signed [w10-1:0] ka568=91;	reg signed [w10-1:0] kb568=-79;	reg signed [w10-1:0] kc568=42;	reg signed [w10-1:0] kd568=-50;	reg signed [w10-1:0] ke568=-11;	reg signed [w10-1:0] kf568=-32;	reg signed [w10-1:0] kg568=34;	reg signed [w10-1:0] kh568=58;	reg signed [w10-1:0] ki568=-105;
reg signed [w10-1:0] ka569=-162;	reg signed [w10-1:0] kb569=-27;	reg signed [w10-1:0] kc569=-60;	reg signed [w10-1:0] kd569=-118;	reg signed [w10-1:0] ke569=10;	reg signed [w10-1:0] kf569=-68;	reg signed [w10-1:0] kg569=120;	reg signed [w10-1:0] kh569=-88;	reg signed [w10-1:0] ki569=-68;
reg signed [w10-1:0] ka570=-109;	reg signed [w10-1:0] kb570=-79;	reg signed [w10-1:0] kc570=88;	reg signed [w10-1:0] kd570=-65;	reg signed [w10-1:0] ke570=-65;	reg signed [w10-1:0] kf570=-76;	reg signed [w10-1:0] kg570=-104;	reg signed [w10-1:0] kh570=61;	reg signed [w10-1:0] ki570=31;
reg signed [w10-1:0] ka571=-25;	reg signed [w10-1:0] kb571=-64;	reg signed [w10-1:0] kc571=75;	reg signed [w10-1:0] kd571=-64;	reg signed [w10-1:0] ke571=90;	reg signed [w10-1:0] kf571=-64;	reg signed [w10-1:0] kg571=-69;	reg signed [w10-1:0] kh571=27;	reg signed [w10-1:0] ki571=-30;
reg signed [w10-1:0] ka572=27;	reg signed [w10-1:0] kb572=-134;	reg signed [w10-1:0] kc572=-19;	reg signed [w10-1:0] kd572=-33;	reg signed [w10-1:0] ke572=99;	reg signed [w10-1:0] kf572=-57;	reg signed [w10-1:0] kg572=78;	reg signed [w10-1:0] kh572=30;	reg signed [w10-1:0] ki572=-36;
reg signed [w10-1:0] ka573=73;	reg signed [w10-1:0] kb573=-54;	reg signed [w10-1:0] kc573=-24;	reg signed [w10-1:0] kd573=-68;	reg signed [w10-1:0] ke573=-57;	reg signed [w10-1:0] kf573=-125;	reg signed [w10-1:0] kg573=74;	reg signed [w10-1:0] kh573=6;	reg signed [w10-1:0] ki573=43;
reg signed [w10-1:0] ka574=-51;	reg signed [w10-1:0] kb574=44;	reg signed [w10-1:0] kc574=-68;	reg signed [w10-1:0] kd574=126;	reg signed [w10-1:0] ke574=127;	reg signed [w10-1:0] kf574=-14;	reg signed [w10-1:0] kg574=-59;	reg signed [w10-1:0] kh574=11;	reg signed [w10-1:0] ki574=77;
reg signed [w10-1:0] ka575=133;	reg signed [w10-1:0] kb575=108;	reg signed [w10-1:0] kc575=-23;	reg signed [w10-1:0] kd575=51;	reg signed [w10-1:0] ke575=-130;	reg signed [w10-1:0] kf575=-47;	reg signed [w10-1:0] kg575=79;	reg signed [w10-1:0] kh575=59;	reg signed [w10-1:0] ki575=-132;
reg signed [w10-1:0] ka576=70;	reg signed [w10-1:0] kb576=0;	reg signed [w10-1:0] kc576=-90;	reg signed [w10-1:0] kd576=23;	reg signed [w10-1:0] ke576=20;	reg signed [w10-1:0] kf576=13;	reg signed [w10-1:0] kg576=-32;	reg signed [w10-1:0] kh576=55;	reg signed [w10-1:0] ki576=20;
reg signed [w10-1:0] ka577=72;	reg signed [w10-1:0] kb577=77;	reg signed [w10-1:0] kc577=44;	reg signed [w10-1:0] kd577=13;	reg signed [w10-1:0] ke577=-7;	reg signed [w10-1:0] kf577=68;	reg signed [w10-1:0] kg577=21;	reg signed [w10-1:0] kh577=76;	reg signed [w10-1:0] ki577=-64;
reg signed [w10-1:0] ka578=112;	reg signed [w10-1:0] kb578=-64;	reg signed [w10-1:0] kc578=107;	reg signed [w10-1:0] kd578=-42;	reg signed [w10-1:0] ke578=-51;	reg signed [w10-1:0] kf578=-69;	reg signed [w10-1:0] kg578=-91;	reg signed [w10-1:0] kh578=49;	reg signed [w10-1:0] ki578=33;
reg signed [w10-1:0] ka579=-113;	reg signed [w10-1:0] kb579=93;	reg signed [w10-1:0] kc579=100;	reg signed [w10-1:0] kd579=-117;	reg signed [w10-1:0] ke579=38;	reg signed [w10-1:0] kf579=133;	reg signed [w10-1:0] kg579=-92;	reg signed [w10-1:0] kh579=-128;	reg signed [w10-1:0] ki579=-14;
reg signed [w10-1:0] ka580=-58;	reg signed [w10-1:0] kb580=60;	reg signed [w10-1:0] kc580=14;	reg signed [w10-1:0] kd580=9;	reg signed [w10-1:0] ke580=112;	reg signed [w10-1:0] kf580=48;	reg signed [w10-1:0] kg580=-62;	reg signed [w10-1:0] kh580=-94;	reg signed [w10-1:0] ki580=-3;
reg signed [w10-1:0] ka581=120;	reg signed [w10-1:0] kb581=10;	reg signed [w10-1:0] kc581=57;	reg signed [w10-1:0] kd581=-92;	reg signed [w10-1:0] ke581=-152;	reg signed [w10-1:0] kf581=-70;	reg signed [w10-1:0] kg581=-102;	reg signed [w10-1:0] kh581=-81;	reg signed [w10-1:0] ki581=42;
reg signed [w10-1:0] ka582=49;	reg signed [w10-1:0] kb582=-46;	reg signed [w10-1:0] kc582=12;	reg signed [w10-1:0] kd582=105;	reg signed [w10-1:0] ke582=44;	reg signed [w10-1:0] kf582=75;	reg signed [w10-1:0] kg582=14;	reg signed [w10-1:0] kh582=54;	reg signed [w10-1:0] ki582=19;
reg signed [w10-1:0] ka583=-93;	reg signed [w10-1:0] kb583=119;	reg signed [w10-1:0] kc583=-69;	reg signed [w10-1:0] kd583=-47;	reg signed [w10-1:0] ke583=-42;	reg signed [w10-1:0] kf583=104;	reg signed [w10-1:0] kg583=68;	reg signed [w10-1:0] kh583=-112;	reg signed [w10-1:0] ki583=77;
reg signed [w10-1:0] ka584=-1;	reg signed [w10-1:0] kb584=-4;	reg signed [w10-1:0] kc584=140;	reg signed [w10-1:0] kd584=43;	reg signed [w10-1:0] ke584=-4;	reg signed [w10-1:0] kf584=-99;	reg signed [w10-1:0] kg584=11;	reg signed [w10-1:0] kh584=143;	reg signed [w10-1:0] ki584=50;
reg signed [w10-1:0] ka585=60;	reg signed [w10-1:0] kb585=13;	reg signed [w10-1:0] kc585=-67;	reg signed [w10-1:0] kd585=-83;	reg signed [w10-1:0] ke585=-111;	reg signed [w10-1:0] kf585=-4;	reg signed [w10-1:0] kg585=-133;	reg signed [w10-1:0] kh585=2;	reg signed [w10-1:0] ki585=32;
reg signed [w10-1:0] ka586=-110;	reg signed [w10-1:0] kb586=35;	reg signed [w10-1:0] kc586=101;	reg signed [w10-1:0] kd586=83;	reg signed [w10-1:0] ke586=-9;	reg signed [w10-1:0] kf586=-76;	reg signed [w10-1:0] kg586=-113;	reg signed [w10-1:0] kh586=32;	reg signed [w10-1:0] ki586=-77;
reg signed [w10-1:0] ka587=-113;	reg signed [w10-1:0] kb587=87;	reg signed [w10-1:0] kc587=43;	reg signed [w10-1:0] kd587=83;	reg signed [w10-1:0] ke587=-84;	reg signed [w10-1:0] kf587=31;	reg signed [w10-1:0] kg587=54;	reg signed [w10-1:0] kh587=-17;	reg signed [w10-1:0] ki587=-49;
reg signed [w10-1:0] ka588=66;	reg signed [w10-1:0] kb588=-87;	reg signed [w10-1:0] kc588=-5;	reg signed [w10-1:0] kd588=-26;	reg signed [w10-1:0] ke588=70;	reg signed [w10-1:0] kf588=42;	reg signed [w10-1:0] kg588=119;	reg signed [w10-1:0] kh588=116;	reg signed [w10-1:0] ki588=70;
reg signed [w10-1:0] ka589=-56;	reg signed [w10-1:0] kb589=132;	reg signed [w10-1:0] kc589=-108;	reg signed [w10-1:0] kd589=76;	reg signed [w10-1:0] ke589=80;	reg signed [w10-1:0] kf589=-118;	reg signed [w10-1:0] kg589=66;	reg signed [w10-1:0] kh589=-1;	reg signed [w10-1:0] ki589=-102;
reg signed [w10-1:0] ka590=48;	reg signed [w10-1:0] kb590=-67;	reg signed [w10-1:0] kc590=34;	reg signed [w10-1:0] kd590=6;	reg signed [w10-1:0] ke590=-101;	reg signed [w10-1:0] kf590=-120;	reg signed [w10-1:0] kg590=64;	reg signed [w10-1:0] kh590=-72;	reg signed [w10-1:0] ki590=101;
reg signed [w10-1:0] ka591=120;	reg signed [w10-1:0] kb591=26;	reg signed [w10-1:0] kc591=-95;	reg signed [w10-1:0] kd591=-25;	reg signed [w10-1:0] ke591=99;	reg signed [w10-1:0] kf591=-20;	reg signed [w10-1:0] kg591=31;	reg signed [w10-1:0] kh591=-6;	reg signed [w10-1:0] ki591=-46;
reg signed [w10-1:0] ka592=66;	reg signed [w10-1:0] kb592=-86;	reg signed [w10-1:0] kc592=-24;	reg signed [w10-1:0] kd592=86;	reg signed [w10-1:0] ke592=-86;	reg signed [w10-1:0] kf592=59;	reg signed [w10-1:0] kg592=36;	reg signed [w10-1:0] kh592=14;	reg signed [w10-1:0] ki592=-19;
reg signed [w10-1:0] ka593=-63;	reg signed [w10-1:0] kb593=-35;	reg signed [w10-1:0] kc593=17;	reg signed [w10-1:0] kd593=-28;	reg signed [w10-1:0] ke593=6;	reg signed [w10-1:0] kf593=-58;	reg signed [w10-1:0] kg593=84;	reg signed [w10-1:0] kh593=-67;	reg signed [w10-1:0] ki593=-64;
reg signed [w10-1:0] ka594=-4;	reg signed [w10-1:0] kb594=108;	reg signed [w10-1:0] kc594=79;	reg signed [w10-1:0] kd594=14;	reg signed [w10-1:0] ke594=63;	reg signed [w10-1:0] kf594=-19;	reg signed [w10-1:0] kg594=22;	reg signed [w10-1:0] kh594=102;	reg signed [w10-1:0] ki594=-58;
reg signed [w10-1:0] ka595=-101;	reg signed [w10-1:0] kb595=1;	reg signed [w10-1:0] kc595=25;	reg signed [w10-1:0] kd595=-49;	reg signed [w10-1:0] ke595=126;	reg signed [w10-1:0] kf595=26;	reg signed [w10-1:0] kg595=-19;	reg signed [w10-1:0] kh595=109;	reg signed [w10-1:0] ki595=-90;
reg signed [w10-1:0] ka596=3;	reg signed [w10-1:0] kb596=-47;	reg signed [w10-1:0] kc596=3;	reg signed [w10-1:0] kd596=87;	reg signed [w10-1:0] ke596=-45;	reg signed [w10-1:0] kf596=-13;	reg signed [w10-1:0] kg596=-95;	reg signed [w10-1:0] kh596=8;	reg signed [w10-1:0] ki596=-47;
reg signed [w10-1:0] ka597=122;	reg signed [w10-1:0] kb597=-83;	reg signed [w10-1:0] kc597=-29;	reg signed [w10-1:0] kd597=72;	reg signed [w10-1:0] ke597=-111;	reg signed [w10-1:0] kf597=-24;	reg signed [w10-1:0] kg597=-138;	reg signed [w10-1:0] kh597=76;	reg signed [w10-1:0] ki597=21;
reg signed [w10-1:0] ka598=-95;	reg signed [w10-1:0] kb598=-20;	reg signed [w10-1:0] kc598=53;	reg signed [w10-1:0] kd598=-132;	reg signed [w10-1:0] ke598=-69;	reg signed [w10-1:0] kf598=62;	reg signed [w10-1:0] kg598=85;	reg signed [w10-1:0] kh598=-53;	reg signed [w10-1:0] ki598=11;
reg signed [w10-1:0] ka599=-7;	reg signed [w10-1:0] kb599=66;	reg signed [w10-1:0] kc599=-96;	reg signed [w10-1:0] kd599=-30;	reg signed [w10-1:0] ke599=-53;	reg signed [w10-1:0] kf599=-1;	reg signed [w10-1:0] kg599=31;	reg signed [w10-1:0] kh599=82;	reg signed [w10-1:0] ki599=-29;
reg signed [w10-1:0] ka600=65;	reg signed [w10-1:0] kb600=-42;	reg signed [w10-1:0] kc600=10;	reg signed [w10-1:0] kd600=-22;	reg signed [w10-1:0] ke600=-62;	reg signed [w10-1:0] kf600=-17;	reg signed [w10-1:0] kg600=96;	reg signed [w10-1:0] kh600=75;	reg signed [w10-1:0] ki600=18;
reg signed [w10-1:0] ka601=22;	reg signed [w10-1:0] kb601=11;	reg signed [w10-1:0] kc601=11;	reg signed [w10-1:0] kd601=-6;	reg signed [w10-1:0] ke601=100;	reg signed [w10-1:0] kf601=110;	reg signed [w10-1:0] kg601=-83;	reg signed [w10-1:0] kh601=84;	reg signed [w10-1:0] ki601=140;
reg signed [w10-1:0] ka602=30;	reg signed [w10-1:0] kb602=74;	reg signed [w10-1:0] kc602=-19;	reg signed [w10-1:0] kd602=58;	reg signed [w10-1:0] ke602=-91;	reg signed [w10-1:0] kf602=-106;	reg signed [w10-1:0] kg602=-16;	reg signed [w10-1:0] kh602=-32;	reg signed [w10-1:0] ki602=95;
reg signed [w10-1:0] ka603=-46;	reg signed [w10-1:0] kb603=-46;	reg signed [w10-1:0] kc603=-126;	reg signed [w10-1:0] kd603=1;	reg signed [w10-1:0] ke603=30;	reg signed [w10-1:0] kf603=-33;	reg signed [w10-1:0] kg603=51;	reg signed [w10-1:0] kh603=17;	reg signed [w10-1:0] ki603=104;
reg signed [w10-1:0] ka604=-12;	reg signed [w10-1:0] kb604=62;	reg signed [w10-1:0] kc604=-71;	reg signed [w10-1:0] kd604=154;	reg signed [w10-1:0] ke604=30;	reg signed [w10-1:0] kf604=62;	reg signed [w10-1:0] kg604=148;	reg signed [w10-1:0] kh604=47;	reg signed [w10-1:0] ki604=-117;
reg signed [w10-1:0] ka605=-108;	reg signed [w10-1:0] kb605=-97;	reg signed [w10-1:0] kc605=-84;	reg signed [w10-1:0] kd605=-84;	reg signed [w10-1:0] ke605=94;	reg signed [w10-1:0] kf605=-93;	reg signed [w10-1:0] kg605=-19;	reg signed [w10-1:0] kh605=8;	reg signed [w10-1:0] ki605=-114;
reg signed [w10-1:0] ka606=-41;	reg signed [w10-1:0] kb606=8;	reg signed [w10-1:0] kc606=-38;	reg signed [w10-1:0] kd606=3;	reg signed [w10-1:0] ke606=9;	reg signed [w10-1:0] kf606=104;	reg signed [w10-1:0] kg606=15;	reg signed [w10-1:0] kh606=-54;	reg signed [w10-1:0] ki606=12;
reg signed [w10-1:0] ka607=-61;	reg signed [w10-1:0] kb607=-68;	reg signed [w10-1:0] kc607=-31;	reg signed [w10-1:0] kd607=9;	reg signed [w10-1:0] ke607=-13;	reg signed [w10-1:0] kf607=10;	reg signed [w10-1:0] kg607=-13;	reg signed [w10-1:0] kh607=85;	reg signed [w10-1:0] ki607=82;
reg signed [w10-1:0] ka608=-115;	reg signed [w10-1:0] kb608=125;	reg signed [w10-1:0] kc608=80;	reg signed [w10-1:0] kd608=-46;	reg signed [w10-1:0] ke608=-30;	reg signed [w10-1:0] kf608=63;	reg signed [w10-1:0] kg608=165;	reg signed [w10-1:0] kh608=-59;	reg signed [w10-1:0] ki608=-56;
reg signed [w10-1:0] ka609=-69;	reg signed [w10-1:0] kb609=105;	reg signed [w10-1:0] kc609=-24;	reg signed [w10-1:0] kd609=-8;	reg signed [w10-1:0] ke609=-45;	reg signed [w10-1:0] kf609=-118;	reg signed [w10-1:0] kg609=-92;	reg signed [w10-1:0] kh609=38;	reg signed [w10-1:0] ki609=-13;
reg signed [w10-1:0] ka610=80;	reg signed [w10-1:0] kb610=159;	reg signed [w10-1:0] kc610=-47;	reg signed [w10-1:0] kd610=149;	reg signed [w10-1:0] ke610=119;	reg signed [w10-1:0] kf610=-111;	reg signed [w10-1:0] kg610=38;	reg signed [w10-1:0] kh610=-32;	reg signed [w10-1:0] ki610=20;
reg signed [w10-1:0] ka611=7;	reg signed [w10-1:0] kb611=24;	reg signed [w10-1:0] kc611=-39;	reg signed [w10-1:0] kd611=58;	reg signed [w10-1:0] ke611=-64;	reg signed [w10-1:0] kf611=84;	reg signed [w10-1:0] kg611=0;	reg signed [w10-1:0] kh611=-86;	reg signed [w10-1:0] ki611=-22;
reg signed [w10-1:0] ka612=66;	reg signed [w10-1:0] kb612=-68;	reg signed [w10-1:0] kc612=26;	reg signed [w10-1:0] kd612=-100;	reg signed [w10-1:0] ke612=-67;	reg signed [w10-1:0] kf612=49;	reg signed [w10-1:0] kg612=6;	reg signed [w10-1:0] kh612=27;	reg signed [w10-1:0] ki612=122;
reg signed [w10-1:0] ka613=-63;	reg signed [w10-1:0] kb613=-50;	reg signed [w10-1:0] kc613=-69;	reg signed [w10-1:0] kd613=-44;	reg signed [w10-1:0] ke613=-55;	reg signed [w10-1:0] kf613=-36;	reg signed [w10-1:0] kg613=54;	reg signed [w10-1:0] kh613=79;	reg signed [w10-1:0] ki613=-110;
reg signed [w10-1:0] ka614=41;	reg signed [w10-1:0] kb614=131;	reg signed [w10-1:0] kc614=-60;	reg signed [w10-1:0] kd614=-27;	reg signed [w10-1:0] ke614=16;	reg signed [w10-1:0] kf614=-91;	reg signed [w10-1:0] kg614=-54;	reg signed [w10-1:0] kh614=-83;	reg signed [w10-1:0] ki614=-35;
reg signed [w10-1:0] ka615=-53;	reg signed [w10-1:0] kb615=107;	reg signed [w10-1:0] kc615=77;	reg signed [w10-1:0] kd615=21;	reg signed [w10-1:0] ke615=-61;	reg signed [w10-1:0] kf615=58;	reg signed [w10-1:0] kg615=-113;	reg signed [w10-1:0] kh615=-90;	reg signed [w10-1:0] ki615=93;
reg signed [w10-1:0] ka616=24;	reg signed [w10-1:0] kb616=98;	reg signed [w10-1:0] kc616=41;	reg signed [w10-1:0] kd616=101;	reg signed [w10-1:0] ke616=47;	reg signed [w10-1:0] kf616=57;	reg signed [w10-1:0] kg616=66;	reg signed [w10-1:0] kh616=57;	reg signed [w10-1:0] ki616=82;
reg signed [w10-1:0] ka617=84;	reg signed [w10-1:0] kb617=127;	reg signed [w10-1:0] kc617=8;	reg signed [w10-1:0] kd617=-53;	reg signed [w10-1:0] ke617=107;	reg signed [w10-1:0] kf617=127;	reg signed [w10-1:0] kg617=-118;	reg signed [w10-1:0] kh617=-89;	reg signed [w10-1:0] ki617=-119;
reg signed [w10-1:0] ka618=28;	reg signed [w10-1:0] kb618=6;	reg signed [w10-1:0] kc618=-14;	reg signed [w10-1:0] kd618=-80;	reg signed [w10-1:0] ke618=-24;	reg signed [w10-1:0] kf618=76;	reg signed [w10-1:0] kg618=63;	reg signed [w10-1:0] kh618=75;	reg signed [w10-1:0] ki618=45;
reg signed [w10-1:0] ka619=-33;	reg signed [w10-1:0] kb619=68;	reg signed [w10-1:0] kc619=-24;	reg signed [w10-1:0] kd619=38;	reg signed [w10-1:0] ke619=114;	reg signed [w10-1:0] kf619=-136;	reg signed [w10-1:0] kg619=48;	reg signed [w10-1:0] kh619=35;	reg signed [w10-1:0] ki619=-103;
reg signed [w10-1:0] ka620=43;	reg signed [w10-1:0] kb620=-13;	reg signed [w10-1:0] kc620=-85;	reg signed [w10-1:0] kd620=85;	reg signed [w10-1:0] ke620=51;	reg signed [w10-1:0] kf620=-138;	reg signed [w10-1:0] kg620=4;	reg signed [w10-1:0] kh620=-133;	reg signed [w10-1:0] ki620=21;
reg signed [w10-1:0] ka621=7;	reg signed [w10-1:0] kb621=-42;	reg signed [w10-1:0] kc621=-95;	reg signed [w10-1:0] kd621=-110;	reg signed [w10-1:0] ke621=-163;	reg signed [w10-1:0] kf621=-11;	reg signed [w10-1:0] kg621=32;	reg signed [w10-1:0] kh621=88;	reg signed [w10-1:0] ki621=49;
reg signed [w10-1:0] ka622=12;	reg signed [w10-1:0] kb622=-60;	reg signed [w10-1:0] kc622=-42;	reg signed [w10-1:0] kd622=-148;	reg signed [w10-1:0] ke622=52;	reg signed [w10-1:0] kf622=125;	reg signed [w10-1:0] kg622=-29;	reg signed [w10-1:0] kh622=112;	reg signed [w10-1:0] ki622=-30;
reg signed [w10-1:0] ka623=-24;	reg signed [w10-1:0] kb623=-2;	reg signed [w10-1:0] kc623=2;	reg signed [w10-1:0] kd623=48;	reg signed [w10-1:0] ke623=-85;	reg signed [w10-1:0] kf623=130;	reg signed [w10-1:0] kg623=-20;	reg signed [w10-1:0] kh623=-41;	reg signed [w10-1:0] ki623=69;
reg signed [w10-1:0] ka624=-12;	reg signed [w10-1:0] kb624=99;	reg signed [w10-1:0] kc624=39;	reg signed [w10-1:0] kd624=-83;	reg signed [w10-1:0] ke624=123;	reg signed [w10-1:0] kf624=8;	reg signed [w10-1:0] kg624=-59;	reg signed [w10-1:0] kh624=4;	reg signed [w10-1:0] ki624=34;
reg signed [w10-1:0] ka625=99;	reg signed [w10-1:0] kb625=0;	reg signed [w10-1:0] kc625=82;	reg signed [w10-1:0] kd625=-112;	reg signed [w10-1:0] ke625=-46;	reg signed [w10-1:0] kf625=-74;	reg signed [w10-1:0] kg625=-14;	reg signed [w10-1:0] kh625=-30;	reg signed [w10-1:0] ki625=-54;
reg signed [w10-1:0] ka626=-91;	reg signed [w10-1:0] kb626=7;	reg signed [w10-1:0] kc626=-65;	reg signed [w10-1:0] kd626=4;	reg signed [w10-1:0] ke626=-36;	reg signed [w10-1:0] kf626=38;	reg signed [w10-1:0] kg626=-95;	reg signed [w10-1:0] kh626=103;	reg signed [w10-1:0] ki626=-5;
reg signed [w10-1:0] ka627=83;	reg signed [w10-1:0] kb627=-109;	reg signed [w10-1:0] kc627=-127;	reg signed [w10-1:0] kd627=-26;	reg signed [w10-1:0] ke627=-26;	reg signed [w10-1:0] kf627=96;	reg signed [w10-1:0] kg627=-38;	reg signed [w10-1:0] kh627=2;	reg signed [w10-1:0] ki627=81;
reg signed [w10-1:0] ka628=61;	reg signed [w10-1:0] kb628=133;	reg signed [w10-1:0] kc628=-85;	reg signed [w10-1:0] kd628=-33;	reg signed [w10-1:0] ke628=36;	reg signed [w10-1:0] kf628=-14;	reg signed [w10-1:0] kg628=61;	reg signed [w10-1:0] kh628=-151;	reg signed [w10-1:0] ki628=28;
reg signed [w10-1:0] ka629=-5;	reg signed [w10-1:0] kb629=-86;	reg signed [w10-1:0] kc629=-30;	reg signed [w10-1:0] kd629=-30;	reg signed [w10-1:0] ke629=6;	reg signed [w10-1:0] kf629=-25;	reg signed [w10-1:0] kg629=-165;	reg signed [w10-1:0] kh629=-37;	reg signed [w10-1:0] ki629=105;
reg signed [w10-1:0] ka630=-67;	reg signed [w10-1:0] kb630=24;	reg signed [w10-1:0] kc630=121;	reg signed [w10-1:0] kd630=-14;	reg signed [w10-1:0] ke630=3;	reg signed [w10-1:0] kf630=2;	reg signed [w10-1:0] kg630=89;	reg signed [w10-1:0] kh630=9;	reg signed [w10-1:0] ki630=-21;
reg signed [w10-1:0] ka631=45;	reg signed [w10-1:0] kb631=-67;	reg signed [w10-1:0] kc631=-116;	reg signed [w10-1:0] kd631=0;	reg signed [w10-1:0] ke631=27;	reg signed [w10-1:0] kf631=-85;	reg signed [w10-1:0] kg631=131;	reg signed [w10-1:0] kh631=-2;	reg signed [w10-1:0] ki631=-119;
reg signed [w10-1:0] ka632=112;	reg signed [w10-1:0] kb632=98;	reg signed [w10-1:0] kc632=-103;	reg signed [w10-1:0] kd632=20;	reg signed [w10-1:0] ke632=155;	reg signed [w10-1:0] kf632=-107;	reg signed [w10-1:0] kg632=117;	reg signed [w10-1:0] kh632=144;	reg signed [w10-1:0] ki632=-8;
reg signed [w10-1:0] ka633=49;	reg signed [w10-1:0] kb633=18;	reg signed [w10-1:0] kc633=150;	reg signed [w10-1:0] kd633=-45;	reg signed [w10-1:0] ke633=-155;	reg signed [w10-1:0] kf633=-68;	reg signed [w10-1:0] kg633=-57;	reg signed [w10-1:0] kh633=-124;	reg signed [w10-1:0] ki633=17;
reg signed [w10-1:0] ka634=-14;	reg signed [w10-1:0] kb634=52;	reg signed [w10-1:0] kc634=-101;	reg signed [w10-1:0] kd634=51;	reg signed [w10-1:0] ke634=115;	reg signed [w10-1:0] kf634=-77;	reg signed [w10-1:0] kg634=91;	reg signed [w10-1:0] kh634=112;	reg signed [w10-1:0] ki634=111;
reg signed [w10-1:0] ka635=-60;	reg signed [w10-1:0] kb635=-63;	reg signed [w10-1:0] kc635=91;	reg signed [w10-1:0] kd635=-79;	reg signed [w10-1:0] ke635=-61;	reg signed [w10-1:0] kf635=63;	reg signed [w10-1:0] kg635=53;	reg signed [w10-1:0] kh635=-11;	reg signed [w10-1:0] ki635=52;
reg signed [w10-1:0] ka636=-51;	reg signed [w10-1:0] kb636=111;	reg signed [w10-1:0] kc636=-125;	reg signed [w10-1:0] kd636=-24;	reg signed [w10-1:0] ke636=110;	reg signed [w10-1:0] kf636=-64;	reg signed [w10-1:0] kg636=96;	reg signed [w10-1:0] kh636=12;	reg signed [w10-1:0] ki636=50;
reg signed [w10-1:0] ka637=116;	reg signed [w10-1:0] kb637=61;	reg signed [w10-1:0] kc637=59;	reg signed [w10-1:0] kd637=58;	reg signed [w10-1:0] ke637=-41;	reg signed [w10-1:0] kf637=73;	reg signed [w10-1:0] kg637=26;	reg signed [w10-1:0] kh637=118;	reg signed [w10-1:0] ki637=26;
reg signed [w10-1:0] ka638=-29;	reg signed [w10-1:0] kb638=-93;	reg signed [w10-1:0] kc638=52;	reg signed [w10-1:0] kd638=-25;	reg signed [w10-1:0] ke638=73;	reg signed [w10-1:0] kf638=-31;	reg signed [w10-1:0] kg638=99;	reg signed [w10-1:0] kh638=-77;	reg signed [w10-1:0] ki638=46;
reg signed [w10-1:0] ka639=-22;	reg signed [w10-1:0] kb639=-43;	reg signed [w10-1:0] kc639=38;	reg signed [w10-1:0] kd639=107;	reg signed [w10-1:0] ke639=-43;	reg signed [w10-1:0] kf639=110;	reg signed [w10-1:0] kg639=-68;	reg signed [w10-1:0] kh639=-89;	reg signed [w10-1:0] ki639=47;
reg signed [w10-1:0] ka640=6;	reg signed [w10-1:0] kb640=138;	reg signed [w10-1:0] kc640=-53;	reg signed [w10-1:0] kd640=-78;	reg signed [w10-1:0] ke640=45;	reg signed [w10-1:0] kf640=-27;	reg signed [w10-1:0] kg640=-83;	reg signed [w10-1:0] kh640=-99;	reg signed [w10-1:0] ki640=-40;
reg signed [w10-1:0] ka641=81;	reg signed [w10-1:0] kb641=-111;	reg signed [w10-1:0] kc641=126;	reg signed [w10-1:0] kd641=11;	reg signed [w10-1:0] ke641=-112;	reg signed [w10-1:0] kf641=137;	reg signed [w10-1:0] kg641=-76;	reg signed [w10-1:0] kh641=94;	reg signed [w10-1:0] ki641=4;
reg signed [w10-1:0] ka642=42;	reg signed [w10-1:0] kb642=-109;	reg signed [w10-1:0] kc642=-75;	reg signed [w10-1:0] kd642=0;	reg signed [w10-1:0] ke642=-118;	reg signed [w10-1:0] kf642=-51;	reg signed [w10-1:0] kg642=12;	reg signed [w10-1:0] kh642=20;	reg signed [w10-1:0] ki642=-49;
reg signed [w10-1:0] ka643=-103;	reg signed [w10-1:0] kb643=-125;	reg signed [w10-1:0] kc643=32;	reg signed [w10-1:0] kd643=100;	reg signed [w10-1:0] ke643=41;	reg signed [w10-1:0] kf643=-98;	reg signed [w10-1:0] kg643=-21;	reg signed [w10-1:0] kh643=-65;	reg signed [w10-1:0] ki643=-74;
reg signed [w10-1:0] ka644=-64;	reg signed [w10-1:0] kb644=87;	reg signed [w10-1:0] kc644=-16;	reg signed [w10-1:0] kd644=-7;	reg signed [w10-1:0] ke644=0;	reg signed [w10-1:0] kf644=89;	reg signed [w10-1:0] kg644=79;	reg signed [w10-1:0] kh644=-69;	reg signed [w10-1:0] ki644=40;
reg signed [w10-1:0] ka645=-70;	reg signed [w10-1:0] kb645=-117;	reg signed [w10-1:0] kc645=27;	reg signed [w10-1:0] kd645=38;	reg signed [w10-1:0] ke645=-139;	reg signed [w10-1:0] kf645=17;	reg signed [w10-1:0] kg645=94;	reg signed [w10-1:0] kh645=-29;	reg signed [w10-1:0] ki645=-81;
reg signed [w10-1:0] ka646=-88;	reg signed [w10-1:0] kb646=-15;	reg signed [w10-1:0] kc646=-94;	reg signed [w10-1:0] kd646=17;	reg signed [w10-1:0] ke646=88;	reg signed [w10-1:0] kf646=58;	reg signed [w10-1:0] kg646=-65;	reg signed [w10-1:0] kh646=38;	reg signed [w10-1:0] ki646=-86;
reg signed [w10-1:0] ka647=-41;	reg signed [w10-1:0] kb647=85;	reg signed [w10-1:0] kc647=32;	reg signed [w10-1:0] kd647=70;	reg signed [w10-1:0] ke647=-35;	reg signed [w10-1:0] kf647=9;	reg signed [w10-1:0] kg647=-60;	reg signed [w10-1:0] kh647=-8;	reg signed [w10-1:0] ki647=31;
reg signed [w10-1:0] ka648=-22;	reg signed [w10-1:0] kb648=-31;	reg signed [w10-1:0] kc648=112;	reg signed [w10-1:0] kd648=57;	reg signed [w10-1:0] ke648=-70;	reg signed [w10-1:0] kf648=99;	reg signed [w10-1:0] kg648=-27;	reg signed [w10-1:0] kh648=-122;	reg signed [w10-1:0] ki648=-29;


reg signed [w7-1:0] delta25=2168;	reg signed [w7-1:0] mu25=591;	reg signed [w7-1:0] beta25=106168;
reg signed [w7-1:0] delta26=1779;	reg signed [w7-1:0] mu26=-289;	reg signed [w7-1:0] beta26=86799;
reg signed [w7-1:0] delta27=1960;	reg signed [w7-1:0] mu27=379;	reg signed [w7-1:0] beta27=51360;
reg signed [w7-1:0] delta28=1409;	reg signed [w7-1:0] mu28=-336;	reg signed [w7-1:0] beta28=44409;
reg signed [w7-1:0] delta29=1089;	reg signed [w7-1:0] mu29=-1232;	reg signed [w7-1:0] beta29=32202;
reg signed [w7-1:0] delta30=1767;	reg signed [w7-1:0] mu30=-2;	reg signed [w7-1:0] beta30=47873;
reg signed [w7-1:0] delta31=1641;	reg signed [w7-1:0] mu31=-483;	reg signed [w7-1:0] beta31=45621;
reg signed [w7-1:0] delta32=1975;	reg signed [w7-1:0] mu32=-18;	reg signed [w7-1:0] beta32=61921;
reg signed [w7-1:0] delta33=1126;	reg signed [w7-1:0] mu33=24;	reg signed [w7-1:0] beta33=17154;
reg signed [w7-1:0] delta34=1419;	reg signed [w7-1:0] mu34=24;	reg signed [w7-1:0] beta34=14135;
reg signed [w7-1:0] delta35=2233;	reg signed [w7-1:0] mu35=88;	reg signed [w7-1:0] beta35=76990;
reg signed [w7-1:0] delta36=2316;	reg signed [w7-1:0] mu36=96;	reg signed [w7-1:0] beta36=41189;
reg signed [w7-1:0] delta37=1853;	reg signed [w7-1:0] mu37=-318;	reg signed [w7-1:0] beta37=67013;
reg signed [w7-1:0] delta38=2086;	reg signed [w7-1:0] mu38=35;	reg signed [w7-1:0] beta38=34000;
reg signed [w7-1:0] delta39=1806;	reg signed [w7-1:0] mu39=264;	reg signed [w7-1:0] beta39=6388;
reg signed [w7-1:0] delta40=1084;	reg signed [w7-1:0] mu40=-1019;	reg signed [w7-1:0] beta40=14091;
reg signed [w13-1:0] delta41=2158;	reg signed [w13-1:0] mu41=-61;	reg signed [w13-1:0] beta41=87182;
reg signed [w13-1:0] delta42=2087;	reg signed [w13-1:0] mu42=315;	reg signed [w13-1:0] beta42=94384;
reg signed [w13-1:0] delta43=1830;	reg signed [w13-1:0] mu43=37;	reg signed [w13-1:0] beta43=74959;
reg signed [w13-1:0] delta44=1958;	reg signed [w13-1:0] mu44=-3;	reg signed [w13-1:0] beta44=50346;
reg signed [w13-1:0] delta45=1070;	reg signed [w13-1:0] mu45=793;	reg signed [w13-1:0] beta45=2265;
reg signed [w13-1:0] delta46=1617;	reg signed [w13-1:0] mu46=-369;	reg signed [w13-1:0] beta46=35900;
reg signed [w13-1:0] delta47=2038;	reg signed [w13-1:0] mu47=646;	reg signed [w13-1:0] beta47=82629;
reg signed [w13-1:0] delta48=1892;	reg signed [w13-1:0] mu48=-605;	reg signed [w13-1:0] beta48=64960;
reg signed [w13-1:0] delta49=1568;	reg signed [w13-1:0] mu49=258;	reg signed [w13-1:0] beta49=-12638;
reg signed [w13-1:0] delta50=1968;	reg signed [w13-1:0] mu50=318;	reg signed [w13-1:0] beta50=71530;
reg signed [w13-1:0] delta51=1898;	reg signed [w13-1:0] mu51=590;	reg signed [w13-1:0] beta51=42418;
reg signed [w13-1:0] delta52=1761;	reg signed [w13-1:0] mu52=-8;	reg signed [w13-1:0] beta52=44697;
reg signed [w13-1:0] delta53=991;	reg signed [w13-1:0] mu53=-150;	reg signed [w13-1:0] beta53=-10393;
reg signed [w13-1:0] delta54=1678;	reg signed [w13-1:0] mu54=280;	reg signed [w13-1:0] beta54=43326;
reg signed [w13-1:0] delta55=1786;	reg signed [w13-1:0] mu55=51;	reg signed [w13-1:0] beta55=35098;
reg signed [w13-1:0] delta56=2126;	reg signed [w13-1:0] mu56=46;	reg signed [w13-1:0] beta56=25869;


reg [5:0]b1=-4;
reg [5:0]b2=25;
reg [5:0]b3=-4;
reg [5:0]b4=-5;
reg [5:0]b5=-9;
reg [5:0]b6=-16;
reg [5:0]b7=-4;
reg [5:0]b8=19;
reg [5:0]b9=-3;
reg [5:0]b10=1;

/* Convolutional layer-1*/
conv1 cir1(clk,rst,inp,oup1,ka1,kb1,kc1,kd1,ke1,kf1,kg1,kh1,ki1,En1);
conv1 cir2(clk,rst,inp,oup2,ka2,kb2,kc2,kd2,ke2,kf2,kg2,kh2,ki2,En2);
conv1 cir3(clk,rst,inp,oup3,ka3,kb3,kc3,kd3,ke3,kf3,kg3,kh3,ki3,En3);
conv1 cir4(clk,rst,inp,oup4,ka4,kb4,kc4,kd4,ke4,kf4,kg4,kh4,ki4,En4);
conv1 cir5(clk,rst,inp,oup5,ka5,kb5,kc5,kd5,ke5,kf5,kg5,kh5,ki5,En5);
conv1 cir6(clk,rst,inp,oup6,ka6,kb6,kc6,kd6,ke6,kf6,kg6,kh6,ki6,En6);
conv1 cir7(clk,rst,inp,oup7,ka7,kb7,kc7,kd7,ke7,kf7,kg7,kh7,ki7,En7);
conv1 cir8(clk,rst,inp,oup8,ka8,kb8,kc8,kd8,ke8,kf8,kg8,kh8,ki8,En8);



/* Batch Normalization-1*/
batch_norma cir10(oup1,delta1,mu1,beta1,ou1);
batch_norma cir11(oup2,delta2,mu2,beta2,ou2);
batch_norma cir12(oup3,delta3,mu3,beta3,ou3);
batch_norma cir13(oup4,delta4,mu4,beta4,ou4);
batch_norma cir14(oup5,delta5,mu5,beta5,ou5);
batch_norma cir15(oup6,delta6,mu6,beta6,ou6);
batch_norma cir16(oup7,delta7,mu7,beta7,ou7);
batch_norma cir17(oup8,delta8,mu8,beta8,ou8);

/* ReLu-1*/
ReLu cir19(ou1,oua1);
ReLu cir20(ou2,oua2);
ReLu cir21(ou3,oua3);
ReLu cir22(ou4,oua4);
ReLu cir23(ou5,oua5);
ReLu cir24(ou6,oua6);
ReLu cir25(ou7,oua7);
ReLu cir26(ou8,oua8);

always@(posedge clk)
begin 
oux1<=oua1;
oux2<=oua2;
oux3<=oua3;
oux4<=oua4;
oux5<=oua5;
oux6<=oua6;
oux7<=oua7;
oux8<=oua8;
if(En1==1'b1)
Ea<=1'b1;
end
/* max pooling-1*/
max_pooling cir28(clk,oux1,~Ea,oub1,E10);
max_pooling cir29(clk,oux2,~Ea,oub2,E11);
max_pooling cir30(clk,oux3,~Ea,oub3,E12);
max_pooling cir31(clk,oux4,~Ea,oub4,E13);
max_pooling cir32(clk,oux5,~Ea,oub5,E14);
max_pooling cir33(clk,oux6,~Ea,oub6,E15);
max_pooling cir34(clk,oux7,~Ea,oub7,E16);
max_pooling cir35(clk,oux8,~Ea,oub8,E17);


assign clk1=E10;
//assign rst1=rst;


always@(posedge E10)
begin
rst1<=1'b0;
ouz1<=oub1;
ouz2<=oub2;
ouz3<=oub3;
ouz4<=oub4;
ouz5<=oub5;
ouz6<=oub6;
ouz7<=oub7;
ouz8<=oub8;
end 

/* Convolutional layer-2*/
conv2 ci1(clk1,rst1,ouz1,oup9,ka9,kb9,kc9,kd9,ke9,kf9,kg9,kh9,ki9,En9);
conv2 ci2(clk1,rst1,ouz2,oup10,ka10,kb10,kc10,kd10,ke10,kf10,kg10,kh10,ki10,En10);
conv2 ci3(clk1,rst1,ouz3,oup11,ka11,kb11,kc11,kd11,ke11,kf11,kg11,kh11,ki11,En11);
conv2 ci4(clk1,rst1,ouz4,oup12,ka12,kb12,kc12,kd12,ke12,kf12,kg12,kh12,ki12,En12);
conv2 ci5(clk1,rst1,ouz5,oup13,ka13,kb13,kc13,kd13,ke13,kf13,kg13,kh13,ki13,En13);
conv2 ci6(clk1,rst1,ouz6,oup14,ka14,kb14,kc14,kd14,ke14,kf14,kg14,kh14,ki14,En14);
conv2 ci7(clk1,rst1,ouz7,oup15,ka15,kb15,kc15,kd15,ke15,kf15,kg15,kh15,ki15,En15);
conv2 ci8(clk1,rst1,ouz8,oup16,ka16,kb16,kc16,kd16,ke16,kf16,kg16,kh16,ki16,En16);

adding_8 co1(oup9,oup10,oup11,oup12,oup13,oup14,oup15, oup16, add1);


conv2 ci9(clk1,rst1,ouz1,oup17,ka17,kb17,kc17,kd17,ke17,kf17,kg17,kh17,ki17,En17);
conv2 ci10(clk1,rst1,ouz2,oup18,ka18,kb18,kc18,kd18,ke18,kf18,kg18,kh18,ki18,En18);
conv2 ci11(clk1,rst1,ouz3,oup19,ka19,kb19,kc19,kd19,ke19,kf19,kg19,kh19,ki19,En19);
conv2 ci12(clk1,rst1,ouz4,oup20,ka20,kb20,kc20,kd20,ke20,kf20,kg20,kh20,ki20,En20);
conv2 ci13(clk1,rst1,ouz5,oup21,ka21,kb21,kc21,kd21,ke21,kf21,kg21,kh21,ki21,En21);
conv2 ci14(clk1,rst1,ouz6,oup22,ka22,kb22,kc22,kd22,ke22,kf22,kg22,kh22,ki22,En22);
conv2 ci15(clk1,rst1,ouz7,oup23,ka23,kb23,kc23,kd23,ke23,kf23,kg23,kh23,ki23,En23);
conv2 ci16(clk1,rst1,ouz8,oup24,ka24,kb24,kc24,kd24,ke24,kf24,kg24,kh24,ki24,En24);

adding_8 co2(oup17,oup18,oup19,oup20,oup21,oup22,oup23, oup24, add2);

conv2 ci17(clk1,rst1,ouz1,oup25,ka25,kb25,kc25,kd25,ke25,kf25,kg25,kh25,ki25,En25);
conv2 ci18(clk1,rst1,ouz2,oup26,ka26,kb26,kc26,kd26,ke26,kf26,kg26,kh26,ki26,En26);
conv2 ci19(clk1,rst1,ouz3,oup27,ka27,kb27,kc27,kd27,ke27,kf27,kg27,kh27,ki27,En27);
conv2 ci20(clk1,rst1,ouz4,oup28,ka28,kb28,kc28,kd28,ke28,kf28,kg28,kh28,ki28,En28);
conv2 ci21(clk1,rst1,ouz5,oup29,ka29,kb29,kc29,kd29,ke29,kf29,kg29,kh29,ki29,En29);
conv2 ci22(clk1,rst1,ouz6,oup30,ka30,kb30,kc30,kd30,ke30,kf30,kg30,kh30,ki30,En30);
conv2 ci23(clk1,rst1,ouz7,oup31,ka31,kb31,kc31,kd31,ke31,kf31,kg31,kh31,ki31,En31);
conv2 ci24(clk1,rst1,ouz8,oup32,ka32,kb32,kc32,kd32,ke32,kf32,kg32,kh32,ki32,En32);

adding_8 co3(oup25,oup26,oup27,oup28,oup29,oup30,oup31, oup32, add3);

conv2 ci25(clk1,rst1,ouz1,oup33,ka33,kb33,kc33,kd33,ke33,kf33,kg33,kh33,ki33,En33);
conv2 ci26(clk1,rst1,ouz2,oup34,ka34,kb34,kc34,kd34,ke34,kf34,kg34,kh34,ki34,En34);
conv2 ci27(clk1,rst1,ouz3,oup35,ka35,kb35,kc35,kd35,ke35,kf35,kg35,kh35,ki35,En35);
conv2 ci28(clk1,rst1,ouz4,oup36,ka36,kb36,kc36,kd36,ke36,kf36,kg36,kh36,ki36,En36);
conv2 ci29(clk1,rst1,ouz5,oup37,ka37,kb37,kc37,kd37,ke37,kf37,kg37,kh37,ki37,En37);
conv2 ci30(clk1,rst1,ouz6,oup38,ka38,kb38,kc38,kd38,ke38,kf38,kg38,kh38,ki38,En38);
conv2 ci31(clk1,rst1,ouz7,oup39,ka39,kb39,kc39,kd39,ke39,kf39,kg39,kh39,ki39,En39);
conv2 ci32(clk1,rst1,ouz8,oup40,ka40,kb40,kc40,kd40,ke40,kf40,kg40,kh40,ki40,En40);

adding_8 co4(oup33,oup34,oup35,oup36,oup37,oup38,oup39, oup40, add4);

conv2 ci33(clk1,rst1,ouz1,oup41,ka41,kb41,kc41,kd41,ke41,kf41,kg41,kh41,ki41,En41);
conv2 ci34(clk1,rst1,ouz2,oup42,ka42,kb42,kc42,kd42,ke42,kf42,kg42,kh42,ki42,En42);
conv2 ci35(clk1,rst1,ouz3,oup43,ka43,kb43,kc43,kd43,ke43,kf43,kg43,kh43,ki43,En43);
conv2 ci36(clk1,rst1,ouz4,oup44,ka44,kb44,kc44,kd44,ke44,kf44,kg44,kh44,ki44,En44);
conv2 ci37(clk1,rst1,ouz5,oup45,ka45,kb45,kc45,kd45,ke45,kf45,kg45,kh45,ki45,En45);
conv2 ci38(clk1,rst1,ouz6,oup46,ka46,kb46,kc46,kd46,ke46,kf46,kg46,kh46,ki46,En46);
conv2 ci39(clk1,rst1,ouz7,oup47,ka47,kb47,kc47,kd47,ke47,kf47,kg47,kh47,ki47,En47);
conv2 ci40(clk1,rst1,ouz8,oup48,ka48,kb48,kc48,kd48,ke48,kf48,kg48,kh48,ki48,En48);

adding_8 co5(oup41,oup42,oup43,oup44,oup45,oup46,oup47, oup48, add5);

conv2 ci41(clk1,rst1,ouz1,oup49,ka49,kb49,kc49,kd49,ke49,kf49,kg49,kh49,ki49,En49);
conv2 ci42(clk1,rst1,ouz2,oup50,ka50,kb50,kc50,kd50,ke50,kf50,kg50,kh50,ki50,En50);
conv2 ci43(clk1,rst1,ouz3,oup51,ka51,kb51,kc51,kd51,ke51,kf51,kg51,kh51,ki51,En51);
conv2 ci44(clk1,rst1,ouz4,oup52,ka52,kb52,kc52,kd52,ke52,kf52,kg52,kh52,ki52,En52);
conv2 ci45(clk1,rst1,ouz5,oup53,ka53,kb53,kc53,kd53,ke53,kf53,kg53,kh53,ki53,En53);
conv2 ci46(clk1,rst1,ouz6,oup54,ka54,kb54,kc54,kd54,ke54,kf54,kg54,kh54,ki54,En54);
conv2 ci47(clk1,rst1,ouz7,oup55,ka55,kb55,kc55,kd55,ke55,kf55,kg55,kh55,ki55,En55);
conv2 ci48(clk1,rst1,ouz8,oup56,ka56,kb56,kc56,kd56,ke56,kf56,kg56,kh56,ki56,En56);

adding_8 co6(oup49,oup50,oup51,oup52,oup53,oup54,oup55, oup56, add6);

conv2 ci49(clk1,rst1,ouz1,oup57,ka57,kb57,kc57,kd57,ke57,kf57,kg57,kh57,ki57,En57);
conv2 ci50(clk1,rst1,ouz2,oup58,ka58,kb58,kc58,kd58,ke58,kf58,kg58,kh58,ki58,En58);
conv2 ci51(clk1,rst1,ouz3,oup59,ka59,kb59,kc59,kd59,ke59,kf59,kg59,kh59,ki59,En59);
conv2 ci52(clk1,rst1,ouz4,oup60,ka60,kb60,kc60,kd60,ke60,kf60,kg60,kh60,ki60,En60);
conv2 ci53(clk1,rst1,ouz5,oup61,ka61,kb61,kc61,kd61,ke61,kf61,kg61,kh61,ki61,En61);
conv2 ci54(clk1,rst1,ouz6,oup62,ka62,kb62,kc62,kd62,ke62,kf62,kg62,kh62,ki62,En62);
conv2 ci55(clk1,rst1,ouz7,oup63,ka63,kb63,kc63,kd63,ke63,kf63,kg63,kh63,ki63,En63);
conv2 ci56(clk1,rst1,ouz8,oup64,ka64,kb64,kc64,kd64,ke64,kf64,kg64,kh64,ki64,En64);

adding_8 co7(oup57,oup58,oup59,oup60,oup61,oup62,oup63, oup64, add7);

conv2 ci57(clk1,rst1,ouz1,oup65,ka65,kb65,kc65,kd65,ke65,kf65,kg65,kh65,ki65,En65);
conv2 ci58(clk1,rst1,ouz2,oup66,ka66,kb66,kc66,kd66,ke66,kf66,kg66,kh66,ki66,En66);
conv2 ci59(clk1,rst1,ouz3,oup67,ka67,kb67,kc67,kd67,ke67,kf67,kg67,kh67,ki67,En67);
conv2 ci60(clk1,rst1,ouz4,oup68,ka68,kb68,kc68,kd68,ke68,kf68,kg68,kh68,ki68,En68);
conv2 ci61(clk1,rst1,ouz5,oup69,ka69,kb69,kc69,kd69,ke69,kf69,kg69,kh69,ki69,En69);
conv2 ci62(clk1,rst1,ouz6,oup70,ka70,kb70,kc70,kd70,ke70,kf70,kg70,kh70,ki70,En70);
conv2 ci63(clk1,rst1,ouz7,oup71,ka71,kb71,kc71,kd71,ke71,kf71,kg71,kh71,ki71,En71);
conv2 ci64(clk1,rst1,ouz8,oup72,ka72,kb72,kc72,kd72,ke72,kf72,kg72,kh72,ki72,En72);

adding_8 co8(oup65,oup66,oup67,oup68,oup69,oup70,oup71, oup72, add8);

conv2 ci65(clk1,rst1,ouz1,oup73,ka73,kb73,kc73,kd73,ke73,kf73,kg73,kh73,ki73,En73);
conv2 ci66(clk1,rst1,ouz2,oup74,ka74,kb74,kc74,kd74,ke74,kf74,kg74,kh74,ki74,En74);
conv2 ci67(clk1,rst1,ouz3,oup75,ka75,kb75,kc75,kd75,ke75,kf75,kg75,kh75,ki75,En75);
conv2 ci68(clk1,rst1,ouz4,oup76,ka76,kb76,kc76,kd76,ke76,kf76,kg76,kh76,ki76,En76);
conv2 ci69(clk1,rst1,ouz5,oup77,ka77,kb77,kc77,kd77,ke77,kf77,kg77,kh77,ki77,En77);
conv2 ci70(clk1,rst1,ouz6,oup78,ka78,kb78,kc78,kd78,ke78,kf78,kg78,kh78,ki78,En78);
conv2 ci71(clk1,rst1,ouz7,oup79,ka79,kb79,kc79,kd79,ke79,kf79,kg79,kh79,ki79,En79);
conv2 ci72(clk1,rst1,ouz8,oup80,ka80,kb80,kc80,kd80,ke80,kf80,kg80,kh80,ki80,En80);

adding_8 co9(oup73,oup74,oup75,oup76,oup77,oup78,oup79, oup80, add9);

conv2 ci73(clk1,rst1,ouz1,oup81,ka81,kb81,kc81,kd81,ke81,kf81,kg81,kh81,ki81,En81);
conv2 ci74(clk1,rst1,ouz2,oup82,ka82,kb82,kc82,kd82,ke82,kf82,kg82,kh82,ki82,En82);
conv2 ci75(clk1,rst1,ouz3,oup83,ka83,kb83,kc83,kd83,ke83,kf83,kg83,kh83,ki83,En83);
conv2 ci76(clk1,rst1,ouz4,oup84,ka84,kb84,kc84,kd84,ke84,kf84,kg84,kh84,ki84,En84);
conv2 ci77(clk1,rst1,ouz5,oup85,ka85,kb85,kc85,kd85,ke85,kf85,kg85,kh85,ki85,En85);
conv2 ci78(clk1,rst1,ouz6,oup86,ka86,kb86,kc86,kd86,ke86,kf86,kg86,kh86,ki86,En86);
conv2 ci79(clk1,rst1,ouz7,oup87,ka87,kb87,kc87,kd87,ke87,kf87,kg87,kh87,ki87,En87);
conv2 ci80(clk1,rst1,ouz8,oup88,ka88,kb88,kc88,kd88,ke88,kf88,kg88,kh88,ki88,En88);

adding_8 co10(oup81,oup82,oup83,oup84,oup85,oup86,oup87, oup88, add10);

conv2 ci81(clk1,rst1,ouz1,oup89,ka89,kb89,kc89,kd89,ke89,kf89,kg89,kh89,ki89,En89);
conv2 ci82(clk1,rst1,ouz2,oup90,ka90,kb90,kc90,kd90,ke90,kf90,kg90,kh90,ki90,En90);
conv2 ci83(clk1,rst1,ouz3,oup91,ka91,kb91,kc91,kd91,ke91,kf91,kg91,kh91,ki91,En91);
conv2 ci84(clk1,rst1,ouz4,oup92,ka92,kb92,kc92,kd92,ke92,kf92,kg92,kh92,ki92,En92);
conv2 ci85(clk1,rst1,ouz5,oup93,ka93,kb93,kc93,kd93,ke93,kf93,kg93,kh93,ki93,En93);
conv2 ci86(clk1,rst1,ouz6,oup94,ka94,kb94,kc94,kd94,ke94,kf94,kg94,kh94,ki94,En94);
conv2 ci87(clk1,rst1,ouz7,oup95,ka95,kb95,kc95,kd95,ke95,kf95,kg95,kh95,ki95,En95);
conv2 ci88(clk1,rst1,ouz8,oup96,ka96,kb96,kc96,kd96,ke96,kf96,kg96,kh96,ki96,En96);

adding_8 co11(oup89,oup90,oup91,oup92,oup93,oup94,oup95, oup96, add11);

conv2 ci89(clk1,rst1,ouz1,oup97,ka97,kb97,kc97,kd97,ke97,kf97,kg97,kh97,ki97,En97);
conv2 ci90(clk1,rst1,ouz2,oup98,ka98,kb98,kc98,kd98,ke98,kf98,kg98,kh98,ki98,En98);
conv2 ci91(clk1,rst1,ouz3,oup99,ka99,kb99,kc99,kd99,ke99,kf99,kg99,kh99,ki99,En99);
conv2 ci92(clk1,rst1,ouz4,oup100,ka100,kb100,kc100,kd100,ke100,kf100,kg100,kh100,ki100,En100);
conv2 ci93(clk1,rst1,ouz5,oup101,ka101,kb101,kc101,kd101,ke101,kf101,kg101,kh101,ki101,En101);
conv2 ci94(clk1,rst1,ouz6,oup102,ka102,kb102,kc102,kd102,ke102,kf102,kg102,kh102,ki102,En102);
conv2 ci95(clk1,rst1,ouz7,oup103,ka103,kb103,kc103,kd103,ke103,kf103,kg103,kh103,ki103,En103);
conv2 ci96(clk1,rst1,ouz8,oup104,ka104,kb104,kc104,kd104,ke104,kf104,kg104,kh104,ki104,En104);

adding_8 co12(oup97,oup98,oup99,oup100,oup101,oup102,oup103, oup104, add12);

conv2 ci97(clk1,rst1,ouz1,oup105,ka105,kb105,kc105,kd105,ke105,kf105,kg105,kh105,ki105,En105);
conv2 ci98(clk1,rst1,ouz2,oup106,ka106,kb106,kc106,kd106,ke106,kf106,kg106,kh106,ki106,En106);
conv2 ci99(clk1,rst1,ouz3,oup107,ka107,kb107,kc107,kd107,ke107,kf107,kg107,kh107,ki107,En107);
conv2 ci100(clk1,rst1,ouz4,oup108,ka108,kb108,kc108,kd108,ke108,kf108,kg108,kh108,ki108,En108);
conv2 ci101(clk1,rst1,ouz5,oup109,ka109,kb109,kc109,kd109,ke109,kf109,kg109,kh109,ki109,En109);
conv2 ci102(clk1,rst1,ouz6,oup110,ka110,kb110,kc110,kd110,ke110,kf110,kg110,kh110,ki110,En110);
conv2 ci103(clk1,rst1,ouz7,oup111,ka111,kb111,kc111,kd111,ke111,kf111,kg111,kh111,ki111,En111);
conv2 ci104(clk1,rst1,ouz8,oup112,ka112,kb112,kc112,kd112,ke112,kf112,kg112,kh112,ki112,En112);

adding_8 co13(oup105,oup106,oup107,oup108,oup109,oup110,oup111, oup112, add13);

conv2 ci105(clk1,rst1,ouz1,oup113,ka113,kb113,kc113,kd113,ke113,kf113,kg113,kh113,ki113,En113);
conv2 ci106(clk1,rst1,ouz2,oup114,ka114,kb114,kc114,kd114,ke114,kf114,kg114,kh114,ki114,En114);
conv2 ci107(clk1,rst1,ouz3,oup115,ka115,kb115,kc115,kd115,ke115,kf115,kg115,kh115,ki115,En115);
conv2 ci108(clk1,rst1,ouz4,oup116,ka116,kb116,kc116,kd116,ke116,kf116,kg116,kh116,ki116,En116);
conv2 ci109(clk1,rst1,ouz5,oup117,ka117,kb117,kc117,kd117,ke117,kf117,kg117,kh117,ki117,En117);
conv2 ci110(clk1,rst1,ouz6,oup118,ka118,kb118,kc118,kd118,ke118,kf118,kg118,kh118,ki118,En118);
conv2 ci111(clk1,rst1,ouz7,oup119,ka119,kb119,kc119,kd119,ke119,kf119,kg119,kh119,ki119,En119);
conv2 ci112(clk1,rst1,ouz8,oup120,ka120,kb120,kc120,kd120,ke120,kf120,kg120,kh120,ki120,En120);

adding_8 co14(oup113,oup114,oup115,oup116,oup117,oup118,oup119, oup120, add14);

conv2 ci113(clk1,rst1,ouz1,oup121,ka121,kb121,kc121,kd121,ke121,kf121,kg121,kh121,ki121,En121);
conv2 ci114(clk1,rst1,ouz2,oup122,ka122,kb122,kc122,kd122,ke122,kf122,kg122,kh122,ki122,En122);
conv2 ci115(clk1,rst1,ouz3,oup123,ka123,kb123,kc123,kd123,ke123,kf123,kg123,kh123,ki123,En123);
conv2 ci116(clk1,rst1,ouz4,oup124,ka124,kb124,kc124,kd124,ke124,kf124,kg124,kh124,ki124,En124);
conv2 ci117(clk1,rst1,ouz5,oup125,ka125,kb125,kc125,kd125,ke125,kf125,kg125,kh125,ki125,En125);
conv2 ci118(clk1,rst1,ouz6,oup126,ka126,kb126,kc126,kd126,ke126,kf126,kg126,kh126,ki126,En126);
conv2 ci119(clk1,rst1,ouz7,oup127,ka127,kb127,kc127,kd127,ke127,kf127,kg127,kh127,ki127,En127);
conv2 ci120(clk1,rst1,ouz8,oup128,ka128,kb128,kc128,kd128,ke128,kf128,kg128,kh128,ki128,En128);

adding_8 co15(oup121,oup122,oup123,oup124,oup125,oup126,oup127, oup128, add15);

conv2 ci121(clk1,rst1,ouz1,oup129,ka129,kb129,kc129,kd129,ke129,kf129,kg129,kh129,ki129,En129);
conv2 ci122(clk1,rst1,ouz2,oup130,ka130,kb130,kc130,kd130,ke130,kf130,kg130,kh130,ki130,En130);
conv2 ci123(clk1,rst1,ouz3,oup131,ka131,kb131,kc131,kd131,ke131,kf131,kg131,kh131,ki131,En131);
conv2 ci124(clk1,rst1,ouz4,oup132,ka132,kb132,kc132,kd132,ke132,kf132,kg132,kh132,ki132,En132);
conv2 ci125(clk1,rst1,ouz5,oup133,ka133,kb133,kc133,kd133,ke133,kf133,kg133,kh133,ki133,En133);
conv2 ci126(clk1,rst1,ouz6,oup134,ka134,kb134,kc134,kd134,ke134,kf134,kg134,kh134,ki134,En134);
conv2 ci127(clk1,rst1,ouz7,oup135,ka135,kb135,kc135,kd135,ke135,kf135,kg135,kh135,ki135,En135);
conv2 ci128(clk1,rst1,ouz8,oup136,ka136,kb136,kc136,kd136,ke136,kf136,kg136,kh136,ki136,En136);

adding_8 co16(oup129,oup130,oup131,oup132,oup133,oup134,oup135, oup136, add16);

/* Batch Normalization layer-2*/
batch_norm2 bn9(add1,delta9,mu9,beta9,bn_ou1);
batch_norm2 bn10(add2,delta10,mu10,beta10,bn_ou2);
batch_norm2 bn11(add3,delta11,mu11,beta11,bn_ou3);
batch_norm2 bn12(add4,delta12,mu12,beta12,bn_ou4);
batch_norm2 bn13(add5,delta13,mu13,beta13,bn_ou5);
batch_norm2 bn14(add6,delta14,mu14,beta14,bn_ou6);
batch_norm2 bn15(add7,delta15,mu15,beta15,bn_ou7);
batch_norm2 bn16(add8,delta16,mu16,beta16,bn_ou8);
batch_norm2 bn17(add9,delta17,mu17,beta17,bn_ou9);
batch_norm2 bn18(add10,delta18,mu18,beta18,bn_ou10);
batch_norm2 bn19(add11,delta19,mu19,beta19,bn_ou11);
batch_norm2 bn20(add12,delta20,mu20,beta20,bn_ou12);
batch_norm2 bn21(add13,delta21,mu21,beta21,bn_ou13);
batch_norm2 bn22(add14,delta22,mu22,beta22,bn_ou14);
batch_norm2 bn23(add15,delta23,mu23,beta23,bn_ou15);
batch_norm2 bn24(add16,delta24,mu24,beta24,bn_ou16);


/* ReLu layer-2*/
ReLu re1(bn_ou1,ro1);
ReLu re2(bn_ou2,ro2);
ReLu re3(bn_ou3,ro3);
ReLu re4(bn_ou4,ro4);
ReLu re5(bn_ou5,ro5);
ReLu re6(bn_ou6,ro6);
ReLu re7(bn_ou7,ro7);
ReLu re8(bn_ou8,ro8);
ReLu re9(bn_ou9,ro9);
ReLu re10(bn_ou10,ro10);
ReLu re11(bn_ou11,ro11);
ReLu re12(bn_ou12,ro12);
ReLu re13(bn_ou13,ro13);
ReLu re14(bn_ou14,ro14);
ReLu re15(bn_ou15,ro15);
ReLu re16(bn_ou16,ro16);

always@(posedge clk1)
begin 
roa1<=ro1;
roa2<=ro2;
roa3<=ro3;
roa4<=ro4;
roa5<=ro5;
roa6<=ro6;
roa7<=ro7;
roa8<=ro8;
roa9<=ro9;
roa10<=ro10;
roa11<=ro11;
roa12<=ro12;
roa13<=ro13;
roa14<=ro14;
roa15<=ro15;
roa16<=ro16;
if(En9==1'b1)
Eb<=1'b1;
end

/* Max pooling-2*/
max_pooling1 mp1(clk1,roa1,~Eb,mp_ou1,enab1);
max_pooling1 mp2(clk1,roa2,~Eb,mp_ou2,enab2);
max_pooling1 mp3(clk1,roa3,~Eb,mp_ou3,enab3);
max_pooling1 mp4(clk1,roa4,~Eb,mp_ou4,enab4);
max_pooling1 mp5(clk1,roa5,~Eb,mp_ou5,enab5);
max_pooling1 mp6(clk1,roa6,~Eb,mp_ou6,enab6);
max_pooling1 mp7(clk1,roa7,~Eb,mp_ou7,enab7);
max_pooling1 mp8(clk1,roa8,~Eb,mp_ou8,enab8);
max_pooling1 mp9(clk1,roa9,~Eb,mp_ou9,enab9);
max_pooling1 mp10(clk1,roa10,~Eb,mp_ou10,enab10);
max_pooling1 mp11(clk1,roa11,~Eb,mp_ou11,enab11);
max_pooling1 mp12(clk1,roa12,~Eb,mp_ou12,enab12);
max_pooling1 mp13(clk1,roa13,~Eb,mp_ou13,enab13);
max_pooling1 mp14(clk1,roa14,~Eb,mp_ou14,enab14);
max_pooling1 mp15(clk1,roa15,~Eb,mp_ou15,enab15);
max_pooling1 mp16(clk1,roa16,~Eb,mp_ou16,enab16);


assign clk3=enab1;
//assign rst1=rst;


always@(posedge enab1)
begin
rst3<=1'b0;
ouf1<=mp_ou1;
ouf2<=mp_ou2;
ouf3<=mp_ou3;
ouf4<=mp_ou4;
ouf5<=mp_ou5;
ouf6<=mp_ou6;
ouf7<=mp_ou7;
ouf8<=mp_ou8;
ouf9<=mp_ou9;
ouf10<=mp_ou10;
ouf11<=mp_ou11;
ouf12<=mp_ou12;
ouf13<=mp_ou13;
ouf14<=mp_ou14;
ouf15<=mp_ou15;
ouf16<=mp_ou16;
end 

/* Convolutional layer-3*/
conv3 ci137(clk3,rst3,ouf1,oud137,ka137,kb137,kc137,kd137,ke137,kf137,kg137,kh137,ki137,En137);
conv3 ci138(clk3,rst3,ouf2,oud138,ka138,kb138,kc138,kd138,ke138,kf138,kg138,kh138,ki138,En138);
conv3 ci139(clk3,rst3,ouf3,oud139,ka139,kb139,kc139,kd139,ke139,kf139,kg139,kh139,ki139,En139);
conv3 ci140(clk3,rst3,ouf4,oud140,ka140,kb140,kc140,kd140,ke140,kf140,kg140,kh140,ki140,En140);
conv3 ci141(clk3,rst3,ouf5,oud141,ka141,kb141,kc141,kd141,ke141,kf141,kg141,kh141,ki141,En141);
conv3 ci142(clk3,rst3,ouf6,oud142,ka142,kb142,kc142,kd142,ke142,kf142,kg142,kh142,ki142,En142);
conv3 ci143(clk3,rst3,ouf7,oud143,ka143,kb143,kc143,kd143,ke143,kf143,kg143,kh143,ki143,En143);
conv3 ci144(clk3,rst3,ouf8,oud144,ka144,kb144,kc144,kd144,ke144,kf144,kg144,kh144,ki144,En144);
conv3 ci145(clk3,rst3,ouf9,oud145,ka145,kb145,kc145,kd145,ke145,kf145,kg145,kh145,ki145,En145);
conv3 ci146(clk3,rst3,ouf10,oud146,ka146,kb146,kc146,kd146,ke146,kf146,kg146,kh146,ki146,En146);
conv3 ci147(clk3,rst3,ouf11,oud147,ka147,kb147,kc147,kd147,ke147,kf147,kg147,kh147,ki147,En147);
conv3 ci148(clk3,rst3,ouf12,oud148,ka148,kb148,kc148,kd148,ke148,kf148,kg148,kh148,ki148,En148);
conv3 ci149(clk3,rst3,ouf13,oud149,ka149,kb149,kc149,kd149,ke149,kf149,kg149,kh149,ki149,En149);
conv3 ci150(clk3,rst3,ouf14,oud150,ka150,kb150,kc150,kd150,ke150,kf150,kg150,kh150,ki150,En150);
conv3 ci151(clk3,rst3,ouf15,oud151,ka151,kb151,kc151,kd151,ke151,kf151,kg151,kh151,ki151,En151);
conv3 ci152(clk3,rst3,ouf16,oud152,ka152,kb152,kc152,kd152,ke152,kf152,kg152,kh152,ki152,En152);
conv3 ci153(clk3,rst3,ouf1,oud153,ka153,kb153,kc153,kd153,ke153,kf153,kg153,kh153,ki153,En153);
conv3 ci154(clk3,rst3,ouf2,oud154,ka154,kb154,kc154,kd154,ke154,kf154,kg154,kh154,ki154,En154);
conv3 ci155(clk3,rst3,ouf3,oud155,ka155,kb155,kc155,kd155,ke155,kf155,kg155,kh155,ki155,En155);
conv3 ci156(clk3,rst3,ouf4,oud156,ka156,kb156,kc156,kd156,ke156,kf156,kg156,kh156,ki156,En156);
conv3 ci157(clk3,rst3,ouf5,oud157,ka157,kb157,kc157,kd157,ke157,kf157,kg157,kh157,ki157,En157);
conv3 ci158(clk3,rst3,ouf6,oud158,ka158,kb158,kc158,kd158,ke158,kf158,kg158,kh158,ki158,En158);
conv3 ci159(clk3,rst3,ouf7,oud159,ka159,kb159,kc159,kd159,ke159,kf159,kg159,kh159,ki159,En159);
conv3 ci160(clk3,rst3,ouf8,oud160,ka160,kb160,kc160,kd160,ke160,kf160,kg160,kh160,ki160,En160);
conv3 ci161(clk3,rst3,ouf9,oud161,ka161,kb161,kc161,kd161,ke161,kf161,kg161,kh161,ki161,En161);
conv3 ci162(clk3,rst3,ouf10,oud162,ka162,kb162,kc162,kd162,ke162,kf162,kg162,kh162,ki162,En162);
conv3 ci163(clk3,rst3,ouf11,oud163,ka163,kb163,kc163,kd163,ke163,kf163,kg163,kh163,ki163,En163);
conv3 ci164(clk3,rst3,ouf12,oud164,ka164,kb164,kc164,kd164,ke164,kf164,kg164,kh164,ki164,En164);
conv3 ci165(clk3,rst3,ouf13,oud165,ka165,kb165,kc165,kd165,ke165,kf165,kg165,kh165,ki165,En165);
conv3 ci166(clk3,rst3,ouf14,oud166,ka166,kb166,kc166,kd166,ke166,kf166,kg166,kh166,ki166,En166);
conv3 ci167(clk3,rst3,ouf15,oud167,ka167,kb167,kc167,kd167,ke167,kf167,kg167,kh167,ki167,En167);
conv3 ci168(clk3,rst3,ouf16,oud168,ka168,kb168,kc168,kd168,ke168,kf168,kg168,kh168,ki168,En168);
conv3 ci169(clk3,rst3,ouf1,oud169,ka169,kb169,kc169,kd169,ke169,kf169,kg169,kh169,ki169,En169);
conv3 ci170(clk3,rst3,ouf2,oud170,ka170,kb170,kc170,kd170,ke170,kf170,kg170,kh170,ki170,En170);
conv3 ci171(clk3,rst3,ouf3,oud171,ka171,kb171,kc171,kd171,ke171,kf171,kg171,kh171,ki171,En171);
conv3 ci172(clk3,rst3,ouf4,oud172,ka172,kb172,kc172,kd172,ke172,kf172,kg172,kh172,ki172,En172);
conv3 ci173(clk3,rst3,ouf5,oud173,ka173,kb173,kc173,kd173,ke173,kf173,kg173,kh173,ki173,En173);
conv3 ci174(clk3,rst3,ouf6,oud174,ka174,kb174,kc174,kd174,ke174,kf174,kg174,kh174,ki174,En174);
conv3 ci175(clk3,rst3,ouf7,oud175,ka175,kb175,kc175,kd175,ke175,kf175,kg175,kh175,ki175,En175);
conv3 ci176(clk3,rst3,ouf8,oud176,ka176,kb176,kc176,kd176,ke176,kf176,kg176,kh176,ki176,En176);
conv3 ci177(clk3,rst3,ouf9,oud177,ka177,kb177,kc177,kd177,ke177,kf177,kg177,kh177,ki177,En177);
conv3 ci178(clk3,rst3,ouf10,oud178,ka178,kb178,kc178,kd178,ke178,kf178,kg178,kh178,ki178,En178);
conv3 ci179(clk3,rst3,ouf11,oud179,ka179,kb179,kc179,kd179,ke179,kf179,kg179,kh179,ki179,En179);
conv3 ci180(clk3,rst3,ouf12,oud180,ka180,kb180,kc180,kd180,ke180,kf180,kg180,kh180,ki180,En180);
conv3 ci181(clk3,rst3,ouf13,oud181,ka181,kb181,kc181,kd181,ke181,kf181,kg181,kh181,ki181,En181);
conv3 ci182(clk3,rst3,ouf14,oud182,ka182,kb182,kc182,kd182,ke182,kf182,kg182,kh182,ki182,En182);
conv3 ci183(clk3,rst3,ouf15,oud183,ka183,kb183,kc183,kd183,ke183,kf183,kg183,kh183,ki183,En183);
conv3 ci184(clk3,rst3,ouf16,oud184,ka184,kb184,kc184,kd184,ke184,kf184,kg184,kh184,ki184,En184);
conv3 ci185(clk3,rst3,ouf1,oud185,ka185,kb185,kc185,kd185,ke185,kf185,kg185,kh185,ki185,En185);
conv3 ci186(clk3,rst3,ouf2,oud186,ka186,kb186,kc186,kd186,ke186,kf186,kg186,kh186,ki186,En186);
conv3 ci187(clk3,rst3,ouf3,oud187,ka187,kb187,kc187,kd187,ke187,kf187,kg187,kh187,ki187,En187);
conv3 ci188(clk3,rst3,ouf4,oud188,ka188,kb188,kc188,kd188,ke188,kf188,kg188,kh188,ki188,En188);
conv3 ci189(clk3,rst3,ouf5,oud189,ka189,kb189,kc189,kd189,ke189,kf189,kg189,kh189,ki189,En189);
conv3 ci190(clk3,rst3,ouf6,oud190,ka190,kb190,kc190,kd190,ke190,kf190,kg190,kh190,ki190,En190);
conv3 ci191(clk3,rst3,ouf7,oud191,ka191,kb191,kc191,kd191,ke191,kf191,kg191,kh191,ki191,En191);
conv3 ci192(clk3,rst3,ouf8,oud192,ka192,kb192,kc192,kd192,ke192,kf192,kg192,kh192,ki192,En192);
conv3 ci193(clk3,rst3,ouf9,oud193,ka193,kb193,kc193,kd193,ke193,kf193,kg193,kh193,ki193,En193);
conv3 ci194(clk3,rst3,ouf10,oud194,ka194,kb194,kc194,kd194,ke194,kf194,kg194,kh194,ki194,En194);
conv3 ci195(clk3,rst3,ouf11,oud195,ka195,kb195,kc195,kd195,ke195,kf195,kg195,kh195,ki195,En195);
conv3 ci196(clk3,rst3,ouf12,oud196,ka196,kb196,kc196,kd196,ke196,kf196,kg196,kh196,ki196,En196);
conv3 ci197(clk3,rst3,ouf13,oud197,ka197,kb197,kc197,kd197,ke197,kf197,kg197,kh197,ki197,En197);
conv3 ci198(clk3,rst3,ouf14,oud198,ka198,kb198,kc198,kd198,ke198,kf198,kg198,kh198,ki198,En198);
conv3 ci199(clk3,rst3,ouf15,oud199,ka199,kb199,kc199,kd199,ke199,kf199,kg199,kh199,ki199,En199);
conv3 ci200(clk3,rst3,ouf16,oud200,ka200,kb200,kc200,kd200,ke200,kf200,kg200,kh200,ki200,En200);
conv3 ci201(clk3,rst3,ouf1,oud201,ka201,kb201,kc201,kd201,ke201,kf201,kg201,kh201,ki201,En201);
conv3 ci202(clk3,rst3,ouf2,oud202,ka202,kb202,kc202,kd202,ke202,kf202,kg202,kh202,ki202,En202);
conv3 ci203(clk3,rst3,ouf3,oud203,ka203,kb203,kc203,kd203,ke203,kf203,kg203,kh203,ki203,En203);
conv3 ci204(clk3,rst3,ouf4,oud204,ka204,kb204,kc204,kd204,ke204,kf204,kg204,kh204,ki204,En204);
conv3 ci205(clk3,rst3,ouf5,oud205,ka205,kb205,kc205,kd205,ke205,kf205,kg205,kh205,ki205,En205);
conv3 ci206(clk3,rst3,ouf6,oud206,ka206,kb206,kc206,kd206,ke206,kf206,kg206,kh206,ki206,En206);
conv3 ci207(clk3,rst3,ouf7,oud207,ka207,kb207,kc207,kd207,ke207,kf207,kg207,kh207,ki207,En207);
conv3 ci208(clk3,rst3,ouf8,oud208,ka208,kb208,kc208,kd208,ke208,kf208,kg208,kh208,ki208,En208);
conv3 ci209(clk3,rst3,ouf9,oud209,ka209,kb209,kc209,kd209,ke209,kf209,kg209,kh209,ki209,En209);
conv3 ci210(clk3,rst3,ouf10,oud210,ka210,kb210,kc210,kd210,ke210,kf210,kg210,kh210,ki210,En210);
conv3 ci211(clk3,rst3,ouf11,oud211,ka211,kb211,kc211,kd211,ke211,kf211,kg211,kh211,ki211,En211);
conv3 ci212(clk3,rst3,ouf12,oud212,ka212,kb212,kc212,kd212,ke212,kf212,kg212,kh212,ki212,En212);
conv3 ci213(clk3,rst3,ouf13,oud213,ka213,kb213,kc213,kd213,ke213,kf213,kg213,kh213,ki213,En213);
conv3 ci214(clk3,rst3,ouf14,oud214,ka214,kb214,kc214,kd214,ke214,kf214,kg214,kh214,ki214,En214);
conv3 ci215(clk3,rst3,ouf15,oud215,ka215,kb215,kc215,kd215,ke215,kf215,kg215,kh215,ki215,En215);
conv3 ci216(clk3,rst3,ouf16,oud216,ka216,kb216,kc216,kd216,ke216,kf216,kg216,kh216,ki216,En216);
conv3 ci217(clk3,rst3,ouf1,oud217,ka217,kb217,kc217,kd217,ke217,kf217,kg217,kh217,ki217,En217);
conv3 ci218(clk3,rst3,ouf2,oud218,ka218,kb218,kc218,kd218,ke218,kf218,kg218,kh218,ki218,En218);
conv3 ci219(clk3,rst3,ouf3,oud219,ka219,kb219,kc219,kd219,ke219,kf219,kg219,kh219,ki219,En219);
conv3 ci220(clk3,rst3,ouf4,oud220,ka220,kb220,kc220,kd220,ke220,kf220,kg220,kh220,ki220,En220);
conv3 ci221(clk3,rst3,ouf5,oud221,ka221,kb221,kc221,kd221,ke221,kf221,kg221,kh221,ki221,En221);
conv3 ci222(clk3,rst3,ouf6,oud222,ka222,kb222,kc222,kd222,ke222,kf222,kg222,kh222,ki222,En222);
conv3 ci223(clk3,rst3,ouf7,oud223,ka223,kb223,kc223,kd223,ke223,kf223,kg223,kh223,ki223,En223);
conv3 ci224(clk3,rst3,ouf8,oud224,ka224,kb224,kc224,kd224,ke224,kf224,kg224,kh224,ki224,En224);
conv3 ci225(clk3,rst3,ouf9,oud225,ka225,kb225,kc225,kd225,ke225,kf225,kg225,kh225,ki225,En225);
conv3 ci226(clk3,rst3,ouf10,oud226,ka226,kb226,kc226,kd226,ke226,kf226,kg226,kh226,ki226,En226);
conv3 ci227(clk3,rst3,ouf11,oud227,ka227,kb227,kc227,kd227,ke227,kf227,kg227,kh227,ki227,En227);
conv3 ci228(clk3,rst3,ouf12,oud228,ka228,kb228,kc228,kd228,ke228,kf228,kg228,kh228,ki228,En228);
conv3 ci229(clk3,rst3,ouf13,oud229,ka229,kb229,kc229,kd229,ke229,kf229,kg229,kh229,ki229,En229);
conv3 ci230(clk3,rst3,ouf14,oud230,ka230,kb230,kc230,kd230,ke230,kf230,kg230,kh230,ki230,En230);
conv3 ci231(clk3,rst3,ouf15,oud231,ka231,kb231,kc231,kd231,ke231,kf231,kg231,kh231,ki231,En231);
conv3 ci232(clk3,rst3,ouf16,oud232,ka232,kb232,kc232,kd232,ke232,kf232,kg232,kh232,ki232,En232);
conv3 ci233(clk3,rst3,ouf1,oud233,ka233,kb233,kc233,kd233,ke233,kf233,kg233,kh233,ki233,En233);
conv3 ci234(clk3,rst3,ouf2,oud234,ka234,kb234,kc234,kd234,ke234,kf234,kg234,kh234,ki234,En234);
conv3 ci235(clk3,rst3,ouf3,oud235,ka235,kb235,kc235,kd235,ke235,kf235,kg235,kh235,ki235,En235);
conv3 ci236(clk3,rst3,ouf4,oud236,ka236,kb236,kc236,kd236,ke236,kf236,kg236,kh236,ki236,En236);
conv3 ci237(clk3,rst3,ouf5,oud237,ka237,kb237,kc237,kd237,ke237,kf237,kg237,kh237,ki237,En237);
conv3 ci238(clk3,rst3,ouf6,oud238,ka238,kb238,kc238,kd238,ke238,kf238,kg238,kh238,ki238,En238);
conv3 ci239(clk3,rst3,ouf7,oud239,ka239,kb239,kc239,kd239,ke239,kf239,kg239,kh239,ki239,En239);
conv3 ci240(clk3,rst3,ouf8,oud240,ka240,kb240,kc240,kd240,ke240,kf240,kg240,kh240,ki240,En240);
conv3 ci241(clk3,rst3,ouf9,oud241,ka241,kb241,kc241,kd241,ke241,kf241,kg241,kh241,ki241,En241);
conv3 ci242(clk3,rst3,ouf10,oud242,ka242,kb242,kc242,kd242,ke242,kf242,kg242,kh242,ki242,En242);
conv3 ci243(clk3,rst3,ouf11,oud243,ka243,kb243,kc243,kd243,ke243,kf243,kg243,kh243,ki243,En243);
conv3 ci244(clk3,rst3,ouf12,oud244,ka244,kb244,kc244,kd244,ke244,kf244,kg244,kh244,ki244,En244);
conv3 ci245(clk3,rst3,ouf13,oud245,ka245,kb245,kc245,kd245,ke245,kf245,kg245,kh245,ki245,En245);
conv3 ci246(clk3,rst3,ouf14,oud246,ka246,kb246,kc246,kd246,ke246,kf246,kg246,kh246,ki246,En246);
conv3 ci247(clk3,rst3,ouf15,oud247,ka247,kb247,kc247,kd247,ke247,kf247,kg247,kh247,ki247,En247);
conv3 ci248(clk3,rst3,ouf16,oud248,ka248,kb248,kc248,kd248,ke248,kf248,kg248,kh248,ki248,En248);
conv3 ci249(clk3,rst3,ouf1,oud249,ka249,kb249,kc249,kd249,ke249,kf249,kg249,kh249,ki249,En249);
conv3 ci250(clk3,rst3,ouf2,oud250,ka250,kb250,kc250,kd250,ke250,kf250,kg250,kh250,ki250,En250);
conv3 ci251(clk3,rst3,ouf3,oud251,ka251,kb251,kc251,kd251,ke251,kf251,kg251,kh251,ki251,En251);
conv3 ci252(clk3,rst3,ouf4,oud252,ka252,kb252,kc252,kd252,ke252,kf252,kg252,kh252,ki252,En252);
conv3 ci253(clk3,rst3,ouf5,oud253,ka253,kb253,kc253,kd253,ke253,kf253,kg253,kh253,ki253,En253);
conv3 ci254(clk3,rst3,ouf6,oud254,ka254,kb254,kc254,kd254,ke254,kf254,kg254,kh254,ki254,En254);
conv3 ci255(clk3,rst3,ouf7,oud255,ka255,kb255,kc255,kd255,ke255,kf255,kg255,kh255,ki255,En255);
conv3 ci256(clk3,rst3,ouf8,oud256,ka256,kb256,kc256,kd256,ke256,kf256,kg256,kh256,ki256,En256);
conv3 ci257(clk3,rst3,ouf9,oud257,ka257,kb257,kc257,kd257,ke257,kf257,kg257,kh257,ki257,En257);
conv3 ci258(clk3,rst3,ouf10,oud258,ka258,kb258,kc258,kd258,ke258,kf258,kg258,kh258,ki258,En258);
conv3 ci259(clk3,rst3,ouf11,oud259,ka259,kb259,kc259,kd259,ke259,kf259,kg259,kh259,ki259,En259);
conv3 ci260(clk3,rst3,ouf12,oud260,ka260,kb260,kc260,kd260,ke260,kf260,kg260,kh260,ki260,En260);
conv3 ci261(clk3,rst3,ouf13,oud261,ka261,kb261,kc261,kd261,ke261,kf261,kg261,kh261,ki261,En261);
conv3 ci262(clk3,rst3,ouf14,oud262,ka262,kb262,kc262,kd262,ke262,kf262,kg262,kh262,ki262,En262);
conv3 ci263(clk3,rst3,ouf15,oud263,ka263,kb263,kc263,kd263,ke263,kf263,kg263,kh263,ki263,En263);
conv3 ci264(clk3,rst3,ouf16,oud264,ka264,kb264,kc264,kd264,ke264,kf264,kg264,kh264,ki264,En264);
conv3 ci265(clk3,rst3,ouf1,oud265,ka265,kb265,kc265,kd265,ke265,kf265,kg265,kh265,ki265,En265);
conv3 ci266(clk3,rst3,ouf2,oud266,ka266,kb266,kc266,kd266,ke266,kf266,kg266,kh266,ki266,En266);
conv3 ci267(clk3,rst3,ouf3,oud267,ka267,kb267,kc267,kd267,ke267,kf267,kg267,kh267,ki267,En267);
conv3 ci268(clk3,rst3,ouf4,oud268,ka268,kb268,kc268,kd268,ke268,kf268,kg268,kh268,ki268,En268);
conv3 ci269(clk3,rst3,ouf5,oud269,ka269,kb269,kc269,kd269,ke269,kf269,kg269,kh269,ki269,En269);
conv3 ci270(clk3,rst3,ouf6,oud270,ka270,kb270,kc270,kd270,ke270,kf270,kg270,kh270,ki270,En270);
conv3 ci271(clk3,rst3,ouf7,oud271,ka271,kb271,kc271,kd271,ke271,kf271,kg271,kh271,ki271,En271);
conv3 ci272(clk3,rst3,ouf8,oud272,ka272,kb272,kc272,kd272,ke272,kf272,kg272,kh272,ki272,En272);
conv3 ci273(clk3,rst3,ouf9,oud273,ka273,kb273,kc273,kd273,ke273,kf273,kg273,kh273,ki273,En273);
conv3 ci274(clk3,rst3,ouf10,oud274,ka274,kb274,kc274,kd274,ke274,kf274,kg274,kh274,ki274,En274);
conv3 ci275(clk3,rst3,ouf11,oud275,ka275,kb275,kc275,kd275,ke275,kf275,kg275,kh275,ki275,En275);
conv3 ci276(clk3,rst3,ouf12,oud276,ka276,kb276,kc276,kd276,ke276,kf276,kg276,kh276,ki276,En276);
conv3 ci277(clk3,rst3,ouf13,oud277,ka277,kb277,kc277,kd277,ke277,kf277,kg277,kh277,ki277,En277);
conv3 ci278(clk3,rst3,ouf14,oud278,ka278,kb278,kc278,kd278,ke278,kf278,kg278,kh278,ki278,En278);
conv3 ci279(clk3,rst3,ouf15,oud279,ka279,kb279,kc279,kd279,ke279,kf279,kg279,kh279,ki279,En279);
conv3 ci280(clk3,rst3,ouf16,oud280,ka280,kb280,kc280,kd280,ke280,kf280,kg280,kh280,ki280,En280);
conv3 ci281(clk3,rst3,ouf1,oud281,ka281,kb281,kc281,kd281,ke281,kf281,kg281,kh281,ki281,En281);
conv3 ci282(clk3,rst3,ouf2,oud282,ka282,kb282,kc282,kd282,ke282,kf282,kg282,kh282,ki282,En282);
conv3 ci283(clk3,rst3,ouf3,oud283,ka283,kb283,kc283,kd283,ke283,kf283,kg283,kh283,ki283,En283);
conv3 ci284(clk3,rst3,ouf4,oud284,ka284,kb284,kc284,kd284,ke284,kf284,kg284,kh284,ki284,En284);
conv3 ci285(clk3,rst3,ouf5,oud285,ka285,kb285,kc285,kd285,ke285,kf285,kg285,kh285,ki285,En285);
conv3 ci286(clk3,rst3,ouf6,oud286,ka286,kb286,kc286,kd286,ke286,kf286,kg286,kh286,ki286,En286);
conv3 ci287(clk3,rst3,ouf7,oud287,ka287,kb287,kc287,kd287,ke287,kf287,kg287,kh287,ki287,En287);
conv3 ci288(clk3,rst3,ouf8,oud288,ka288,kb288,kc288,kd288,ke288,kf288,kg288,kh288,ki288,En288);
conv3 ci289(clk3,rst3,ouf9,oud289,ka289,kb289,kc289,kd289,ke289,kf289,kg289,kh289,ki289,En289);
conv3 ci290(clk3,rst3,ouf10,oud290,ka290,kb290,kc290,kd290,ke290,kf290,kg290,kh290,ki290,En290);
conv3 ci291(clk3,rst3,ouf11,oud291,ka291,kb291,kc291,kd291,ke291,kf291,kg291,kh291,ki291,En291);
conv3 ci292(clk3,rst3,ouf12,oud292,ka292,kb292,kc292,kd292,ke292,kf292,kg292,kh292,ki292,En292);
conv3 ci293(clk3,rst3,ouf13,oud293,ka293,kb293,kc293,kd293,ke293,kf293,kg293,kh293,ki293,En293);
conv3 ci294(clk3,rst3,ouf14,oud294,ka294,kb294,kc294,kd294,ke294,kf294,kg294,kh294,ki294,En294);
conv3 ci295(clk3,rst3,ouf15,oud295,ka295,kb295,kc295,kd295,ke295,kf295,kg295,kh295,ki295,En295);
conv3 ci296(clk3,rst3,ouf16,oud296,ka296,kb296,kc296,kd296,ke296,kf296,kg296,kh296,ki296,En296);
conv3 ci297(clk3,rst3,ouf1,oud297,ka297,kb297,kc297,kd297,ke297,kf297,kg297,kh297,ki297,En297);
conv3 ci298(clk3,rst3,ouf2,oud298,ka298,kb298,kc298,kd298,ke298,kf298,kg298,kh298,ki298,En298);
conv3 ci299(clk3,rst3,ouf3,oud299,ka299,kb299,kc299,kd299,ke299,kf299,kg299,kh299,ki299,En299);
conv3 ci300(clk3,rst3,ouf4,oud300,ka300,kb300,kc300,kd300,ke300,kf300,kg300,kh300,ki300,En300);
conv3 ci301(clk3,rst3,ouf5,oud301,ka301,kb301,kc301,kd301,ke301,kf301,kg301,kh301,ki301,En301);
conv3 ci302(clk3,rst3,ouf6,oud302,ka302,kb302,kc302,kd302,ke302,kf302,kg302,kh302,ki302,En302);
conv3 ci303(clk3,rst3,ouf7,oud303,ka303,kb303,kc303,kd303,ke303,kf303,kg303,kh303,ki303,En303);
conv3 ci304(clk3,rst3,ouf8,oud304,ka304,kb304,kc304,kd304,ke304,kf304,kg304,kh304,ki304,En304);
conv3 ci305(clk3,rst3,ouf9,oud305,ka305,kb305,kc305,kd305,ke305,kf305,kg305,kh305,ki305,En305);
conv3 ci306(clk3,rst3,ouf10,oud306,ka306,kb306,kc306,kd306,ke306,kf306,kg306,kh306,ki306,En306);
conv3 ci307(clk3,rst3,ouf11,oud307,ka307,kb307,kc307,kd307,ke307,kf307,kg307,kh307,ki307,En307);
conv3 ci308(clk3,rst3,ouf12,oud308,ka308,kb308,kc308,kd308,ke308,kf308,kg308,kh308,ki308,En308);
conv3 ci309(clk3,rst3,ouf13,oud309,ka309,kb309,kc309,kd309,ke309,kf309,kg309,kh309,ki309,En309);
conv3 ci310(clk3,rst3,ouf14,oud310,ka310,kb310,kc310,kd310,ke310,kf310,kg310,kh310,ki310,En310);
conv3 ci311(clk3,rst3,ouf15,oud311,ka311,kb311,kc311,kd311,ke311,kf311,kg311,kh311,ki311,En311);
conv3 ci312(clk3,rst3,ouf16,oud312,ka312,kb312,kc312,kd312,ke312,kf312,kg312,kh312,ki312,En312);
conv3 ci313(clk3,rst3,ouf1,oud313,ka313,kb313,kc313,kd313,ke313,kf313,kg313,kh313,ki313,En313);
conv3 ci314(clk3,rst3,ouf2,oud314,ka314,kb314,kc314,kd314,ke314,kf314,kg314,kh314,ki314,En314);
conv3 ci315(clk3,rst3,ouf3,oud315,ka315,kb315,kc315,kd315,ke315,kf315,kg315,kh315,ki315,En315);
conv3 ci316(clk3,rst3,ouf4,oud316,ka316,kb316,kc316,kd316,ke316,kf316,kg316,kh316,ki316,En316);
conv3 ci317(clk3,rst3,ouf5,oud317,ka317,kb317,kc317,kd317,ke317,kf317,kg317,kh317,ki317,En317);
conv3 ci318(clk3,rst3,ouf6,oud318,ka318,kb318,kc318,kd318,ke318,kf318,kg318,kh318,ki318,En318);
conv3 ci319(clk3,rst3,ouf7,oud319,ka319,kb319,kc319,kd319,ke319,kf319,kg319,kh319,ki319,En319);
conv3 ci320(clk3,rst3,ouf8,oud320,ka320,kb320,kc320,kd320,ke320,kf320,kg320,kh320,ki320,En320);
conv3 ci321(clk3,rst3,ouf9,oud321,ka321,kb321,kc321,kd321,ke321,kf321,kg321,kh321,ki321,En321);
conv3 ci322(clk3,rst3,ouf10,oud322,ka322,kb322,kc322,kd322,ke322,kf322,kg322,kh322,ki322,En322);
conv3 ci323(clk3,rst3,ouf11,oud323,ka323,kb323,kc323,kd323,ke323,kf323,kg323,kh323,ki323,En323);
conv3 ci324(clk3,rst3,ouf12,oud324,ka324,kb324,kc324,kd324,ke324,kf324,kg324,kh324,ki324,En324);
conv3 ci325(clk3,rst3,ouf13,oud325,ka325,kb325,kc325,kd325,ke325,kf325,kg325,kh325,ki325,En325);
conv3 ci326(clk3,rst3,ouf14,oud326,ka326,kb326,kc326,kd326,ke326,kf326,kg326,kh326,ki326,En326);
conv3 ci327(clk3,rst3,ouf15,oud327,ka327,kb327,kc327,kd327,ke327,kf327,kg327,kh327,ki327,En327);
conv3 ci328(clk3,rst3,ouf16,oud328,ka328,kb328,kc328,kd328,ke328,kf328,kg328,kh328,ki328,En328);
conv3 ci329(clk3,rst3,ouf1,oud329,ka329,kb329,kc329,kd329,ke329,kf329,kg329,kh329,ki329,En329);
conv3 ci330(clk3,rst3,ouf2,oud330,ka330,kb330,kc330,kd330,ke330,kf330,kg330,kh330,ki330,En330);
conv3 ci331(clk3,rst3,ouf3,oud331,ka331,kb331,kc331,kd331,ke331,kf331,kg331,kh331,ki331,En331);
conv3 ci332(clk3,rst3,ouf4,oud332,ka332,kb332,kc332,kd332,ke332,kf332,kg332,kh332,ki332,En332);
conv3 ci333(clk3,rst3,ouf5,oud333,ka333,kb333,kc333,kd333,ke333,kf333,kg333,kh333,ki333,En333);
conv3 ci334(clk3,rst3,ouf6,oud334,ka334,kb334,kc334,kd334,ke334,kf334,kg334,kh334,ki334,En334);
conv3 ci335(clk3,rst3,ouf7,oud335,ka335,kb335,kc335,kd335,ke335,kf335,kg335,kh335,ki335,En335);
conv3 ci336(clk3,rst3,ouf8,oud336,ka336,kb336,kc336,kd336,ke336,kf336,kg336,kh336,ki336,En336);
conv3 ci337(clk3,rst3,ouf9,oud337,ka337,kb337,kc337,kd337,ke337,kf337,kg337,kh337,ki337,En337);
conv3 ci338(clk3,rst3,ouf10,oud338,ka338,kb338,kc338,kd338,ke338,kf338,kg338,kh338,ki338,En338);
conv3 ci339(clk3,rst3,ouf11,oud339,ka339,kb339,kc339,kd339,ke339,kf339,kg339,kh339,ki339,En339);
conv3 ci340(clk3,rst3,ouf12,oud340,ka340,kb340,kc340,kd340,ke340,kf340,kg340,kh340,ki340,En340);
conv3 ci341(clk3,rst3,ouf13,oud341,ka341,kb341,kc341,kd341,ke341,kf341,kg341,kh341,ki341,En341);
conv3 ci342(clk3,rst3,ouf14,oud342,ka342,kb342,kc342,kd342,ke342,kf342,kg342,kh342,ki342,En342);
conv3 ci343(clk3,rst3,ouf15,oud343,ka343,kb343,kc343,kd343,ke343,kf343,kg343,kh343,ki343,En343);
conv3 ci344(clk3,rst3,ouf16,oud344,ka344,kb344,kc344,kd344,ke344,kf344,kg344,kh344,ki344,En344);
conv3 ci345(clk3,rst3,ouf1,oud345,ka345,kb345,kc345,kd345,ke345,kf345,kg345,kh345,ki345,En345);
conv3 ci346(clk3,rst3,ouf2,oud346,ka346,kb346,kc346,kd346,ke346,kf346,kg346,kh346,ki346,En346);
conv3 ci347(clk3,rst3,ouf3,oud347,ka347,kb347,kc347,kd347,ke347,kf347,kg347,kh347,ki347,En347);
conv3 ci348(clk3,rst3,ouf4,oud348,ka348,kb348,kc348,kd348,ke348,kf348,kg348,kh348,ki348,En348);
conv3 ci349(clk3,rst3,ouf5,oud349,ka349,kb349,kc349,kd349,ke349,kf349,kg349,kh349,ki349,En349);
conv3 ci350(clk3,rst3,ouf6,oud350,ka350,kb350,kc350,kd350,ke350,kf350,kg350,kh350,ki350,En350);
conv3 ci351(clk3,rst3,ouf7,oud351,ka351,kb351,kc351,kd351,ke351,kf351,kg351,kh351,ki351,En351);
conv3 ci352(clk3,rst3,ouf8,oud352,ka352,kb352,kc352,kd352,ke352,kf352,kg352,kh352,ki352,En352);
conv3 ci353(clk3,rst3,ouf9,oud353,ka353,kb353,kc353,kd353,ke353,kf353,kg353,kh353,ki353,En353);
conv3 ci354(clk3,rst3,ouf10,oud354,ka354,kb354,kc354,kd354,ke354,kf354,kg354,kh354,ki354,En354);
conv3 ci355(clk3,rst3,ouf11,oud355,ka355,kb355,kc355,kd355,ke355,kf355,kg355,kh355,ki355,En355);
conv3 ci356(clk3,rst3,ouf12,oud356,ka356,kb356,kc356,kd356,ke356,kf356,kg356,kh356,ki356,En356);
conv3 ci357(clk3,rst3,ouf13,oud357,ka357,kb357,kc357,kd357,ke357,kf357,kg357,kh357,ki357,En357);
conv3 ci358(clk3,rst3,ouf14,oud358,ka358,kb358,kc358,kd358,ke358,kf358,kg358,kh358,ki358,En358);
conv3 ci359(clk3,rst3,ouf15,oud359,ka359,kb359,kc359,kd359,ke359,kf359,kg359,kh359,ki359,En359);
conv3 ci360(clk3,rst3,ouf16,oud360,ka360,kb360,kc360,kd360,ke360,kf360,kg360,kh360,ki360,En360);
conv3 ci361(clk3,rst3,ouf1,oud361,ka361,kb361,kc361,kd361,ke361,kf361,kg361,kh361,ki361,En361);
conv3 ci362(clk3,rst3,ouf2,oud362,ka362,kb362,kc362,kd362,ke362,kf362,kg362,kh362,ki362,En362);
conv3 ci363(clk3,rst3,ouf3,oud363,ka363,kb363,kc363,kd363,ke363,kf363,kg363,kh363,ki363,En363);
conv3 ci364(clk3,rst3,ouf4,oud364,ka364,kb364,kc364,kd364,ke364,kf364,kg364,kh364,ki364,En364);
conv3 ci365(clk3,rst3,ouf5,oud365,ka365,kb365,kc365,kd365,ke365,kf365,kg365,kh365,ki365,En365);
conv3 ci366(clk3,rst3,ouf6,oud366,ka366,kb366,kc366,kd366,ke366,kf366,kg366,kh366,ki366,En366);
conv3 ci367(clk3,rst3,ouf7,oud367,ka367,kb367,kc367,kd367,ke367,kf367,kg367,kh367,ki367,En367);
conv3 ci368(clk3,rst3,ouf8,oud368,ka368,kb368,kc368,kd368,ke368,kf368,kg368,kh368,ki368,En368);
conv3 ci369(clk3,rst3,ouf9,oud369,ka369,kb369,kc369,kd369,ke369,kf369,kg369,kh369,ki369,En369);
conv3 ci370(clk3,rst3,ouf10,oud370,ka370,kb370,kc370,kd370,ke370,kf370,kg370,kh370,ki370,En370);
conv3 ci371(clk3,rst3,ouf11,oud371,ka371,kb371,kc371,kd371,ke371,kf371,kg371,kh371,ki371,En371);
conv3 ci372(clk3,rst3,ouf12,oud372,ka372,kb372,kc372,kd372,ke372,kf372,kg372,kh372,ki372,En372);
conv3 ci373(clk3,rst3,ouf13,oud373,ka373,kb373,kc373,kd373,ke373,kf373,kg373,kh373,ki373,En373);
conv3 ci374(clk3,rst3,ouf14,oud374,ka374,kb374,kc374,kd374,ke374,kf374,kg374,kh374,ki374,En374);
conv3 ci375(clk3,rst3,ouf15,oud375,ka375,kb375,kc375,kd375,ke375,kf375,kg375,kh375,ki375,En375);
conv3 ci376(clk3,rst3,ouf16,oud376,ka376,kb376,kc376,kd376,ke376,kf376,kg376,kh376,ki376,En376);
conv3 ci377(clk3,rst3,ouf1,oud377,ka377,kb377,kc377,kd377,ke377,kf377,kg377,kh377,ki377,En377);
conv3 ci378(clk3,rst3,ouf2,oud378,ka378,kb378,kc378,kd378,ke378,kf378,kg378,kh378,ki378,En378);
conv3 ci379(clk3,rst3,ouf3,oud379,ka379,kb379,kc379,kd379,ke379,kf379,kg379,kh379,ki379,En379);
conv3 ci380(clk3,rst3,ouf4,oud380,ka380,kb380,kc380,kd380,ke380,kf380,kg380,kh380,ki380,En380);
conv3 ci381(clk3,rst3,ouf5,oud381,ka381,kb381,kc381,kd381,ke381,kf381,kg381,kh381,ki381,En381);
conv3 ci382(clk3,rst3,ouf6,oud382,ka382,kb382,kc382,kd382,ke382,kf382,kg382,kh382,ki382,En382);
conv3 ci383(clk3,rst3,ouf7,oud383,ka383,kb383,kc383,kd383,ke383,kf383,kg383,kh383,ki383,En383);
conv3 ci384(clk3,rst3,ouf8,oud384,ka384,kb384,kc384,kd384,ke384,kf384,kg384,kh384,ki384,En384);
conv3 ci385(clk3,rst3,ouf9,oud385,ka385,kb385,kc385,kd385,ke385,kf385,kg385,kh385,ki385,En385);
conv3 ci386(clk3,rst3,ouf10,oud386,ka386,kb386,kc386,kd386,ke386,kf386,kg386,kh386,ki386,En386);
conv3 ci387(clk3,rst3,ouf11,oud387,ka387,kb387,kc387,kd387,ke387,kf387,kg387,kh387,ki387,En387);
conv3 ci388(clk3,rst3,ouf12,oud388,ka388,kb388,kc388,kd388,ke388,kf388,kg388,kh388,ki388,En388);
conv3 ci389(clk3,rst3,ouf13,oud389,ka389,kb389,kc389,kd389,ke389,kf389,kg389,kh389,ki389,En389);
conv3 ci390(clk3,rst3,ouf14,oud390,ka390,kb390,kc390,kd390,ke390,kf390,kg390,kh390,ki390,En390);
conv3 ci391(clk3,rst3,ouf15,oud391,ka391,kb391,kc391,kd391,ke391,kf391,kg391,kh391,ki391,En391);
conv3 ci392(clk3,rst3,ouf16,oud392,ka392,kb392,kc392,kd392,ke392,kf392,kg392,kh392,ki392,En392);
conv3 ci393(clk3,rst3,ouf1,oud393,ka393,kb393,kc393,kd393,ke393,kf393,kg393,kh393,ki393,En393);
conv3 ci394(clk3,rst3,ouf2,oud394,ka394,kb394,kc394,kd394,ke394,kf394,kg394,kh394,ki394,En394);
conv3 ci395(clk3,rst3,ouf3,oud395,ka395,kb395,kc395,kd395,ke395,kf395,kg395,kh395,ki395,En395);
conv3 ci396(clk3,rst3,ouf4,oud396,ka396,kb396,kc396,kd396,ke396,kf396,kg396,kh396,ki396,En396);
conv3 ci397(clk3,rst3,ouf5,oud397,ka397,kb397,kc397,kd397,ke397,kf397,kg397,kh397,ki397,En397);
conv3 ci398(clk3,rst3,ouf6,oud398,ka398,kb398,kc398,kd398,ke398,kf398,kg398,kh398,ki398,En398);
conv3 ci399(clk3,rst3,ouf7,oud399,ka399,kb399,kc399,kd399,ke399,kf399,kg399,kh399,ki399,En399);
conv3 ci400(clk3,rst3,ouf8,oud400,ka400,kb400,kc400,kd400,ke400,kf400,kg400,kh400,ki400,En400);
conv3 ci401(clk3,rst3,ouf9,oud401,ka401,kb401,kc401,kd401,ke401,kf401,kg401,kh401,ki401,En401);
conv3 ci402(clk3,rst3,ouf10,oud402,ka402,kb402,kc402,kd402,ke402,kf402,kg402,kh402,ki402,En402);
conv3 ci403(clk3,rst3,ouf11,oud403,ka403,kb403,kc403,kd403,ke403,kf403,kg403,kh403,ki403,En403);
conv3 ci404(clk3,rst3,ouf12,oud404,ka404,kb404,kc404,kd404,ke404,kf404,kg404,kh404,ki404,En404);
conv3 ci405(clk3,rst3,ouf13,oud405,ka405,kb405,kc405,kd405,ke405,kf405,kg405,kh405,ki405,En405);
conv3 ci406(clk3,rst3,ouf14,oud406,ka406,kb406,kc406,kd406,ke406,kf406,kg406,kh406,ki406,En406);
conv3 ci407(clk3,rst3,ouf15,oud407,ka407,kb407,kc407,kd407,ke407,kf407,kg407,kh407,ki407,En407);
conv3 ci408(clk3,rst3,ouf16,oud408,ka408,kb408,kc408,kd408,ke408,kf408,kg408,kh408,ki408,En408);
conv3 ci409(clk3,rst3,ouf1,oud409,ka409,kb409,kc409,kd409,ke409,kf409,kg409,kh409,ki409,En409);
conv3 ci410(clk3,rst3,ouf2,oud410,ka410,kb410,kc410,kd410,ke410,kf410,kg410,kh410,ki410,En410);
conv3 ci411(clk3,rst3,ouf3,oud411,ka411,kb411,kc411,kd411,ke411,kf411,kg411,kh411,ki411,En411);
conv3 ci412(clk3,rst3,ouf4,oud412,ka412,kb412,kc412,kd412,ke412,kf412,kg412,kh412,ki412,En412);
conv3 ci413(clk3,rst3,ouf5,oud413,ka413,kb413,kc413,kd413,ke413,kf413,kg413,kh413,ki413,En413);
conv3 ci414(clk3,rst3,ouf6,oud414,ka414,kb414,kc414,kd414,ke414,kf414,kg414,kh414,ki414,En414);
conv3 ci415(clk3,rst3,ouf7,oud415,ka415,kb415,kc415,kd415,ke415,kf415,kg415,kh415,ki415,En415);
conv3 ci416(clk3,rst3,ouf8,oud416,ka416,kb416,kc416,kd416,ke416,kf416,kg416,kh416,ki416,En416);
conv3 ci417(clk3,rst3,ouf9,oud417,ka417,kb417,kc417,kd417,ke417,kf417,kg417,kh417,ki417,En417);
conv3 ci418(clk3,rst3,ouf10,oud418,ka418,kb418,kc418,kd418,ke418,kf418,kg418,kh418,ki418,En418);
conv3 ci419(clk3,rst3,ouf11,oud419,ka419,kb419,kc419,kd419,ke419,kf419,kg419,kh419,ki419,En419);
conv3 ci420(clk3,rst3,ouf12,oud420,ka420,kb420,kc420,kd420,ke420,kf420,kg420,kh420,ki420,En420);
conv3 ci421(clk3,rst3,ouf13,oud421,ka421,kb421,kc421,kd421,ke421,kf421,kg421,kh421,ki421,En421);
conv3 ci422(clk3,rst3,ouf14,oud422,ka422,kb422,kc422,kd422,ke422,kf422,kg422,kh422,ki422,En422);
conv3 ci423(clk3,rst3,ouf15,oud423,ka423,kb423,kc423,kd423,ke423,kf423,kg423,kh423,ki423,En423);
conv3 ci424(clk3,rst3,ouf16,oud424,ka424,kb424,kc424,kd424,ke424,kf424,kg424,kh424,ki424,En424);
conv3 ci425(clk3,rst3,ouf1,oud425,ka425,kb425,kc425,kd425,ke425,kf425,kg425,kh425,ki425,En425);
conv3 ci426(clk3,rst3,ouf2,oud426,ka426,kb426,kc426,kd426,ke426,kf426,kg426,kh426,ki426,En426);
conv3 ci427(clk3,rst3,ouf3,oud427,ka427,kb427,kc427,kd427,ke427,kf427,kg427,kh427,ki427,En427);
conv3 ci428(clk3,rst3,ouf4,oud428,ka428,kb428,kc428,kd428,ke428,kf428,kg428,kh428,ki428,En428);
conv3 ci429(clk3,rst3,ouf5,oud429,ka429,kb429,kc429,kd429,ke429,kf429,kg429,kh429,ki429,En429);
conv3 ci430(clk3,rst3,ouf6,oud430,ka430,kb430,kc430,kd430,ke430,kf430,kg430,kh430,ki430,En430);
conv3 ci431(clk3,rst3,ouf7,oud431,ka431,kb431,kc431,kd431,ke431,kf431,kg431,kh431,ki431,En431);
conv3 ci432(clk3,rst3,ouf8,oud432,ka432,kb432,kc432,kd432,ke432,kf432,kg432,kh432,ki432,En432);
conv3 ci433(clk3,rst3,ouf9,oud433,ka433,kb433,kc433,kd433,ke433,kf433,kg433,kh433,ki433,En433);
conv3 ci434(clk3,rst3,ouf10,oud434,ka434,kb434,kc434,kd434,ke434,kf434,kg434,kh434,ki434,En434);
conv3 ci435(clk3,rst3,ouf11,oud435,ka435,kb435,kc435,kd435,ke435,kf435,kg435,kh435,ki435,En435);
conv3 ci436(clk3,rst3,ouf12,oud436,ka436,kb436,kc436,kd436,ke436,kf436,kg436,kh436,ki436,En436);
conv3 ci437(clk3,rst3,ouf13,oud437,ka437,kb437,kc437,kd437,ke437,kf437,kg437,kh437,ki437,En437);
conv3 ci438(clk3,rst3,ouf14,oud438,ka438,kb438,kc438,kd438,ke438,kf438,kg438,kh438,ki438,En438);
conv3 ci439(clk3,rst3,ouf15,oud439,ka439,kb439,kc439,kd439,ke439,kf439,kg439,kh439,ki439,En439);
conv3 ci440(clk3,rst3,ouf16,oud440,ka440,kb440,kc440,kd440,ke440,kf440,kg440,kh440,ki440,En440);
conv3 ci441(clk3,rst3,ouf1,oud441,ka441,kb441,kc441,kd441,ke441,kf441,kg441,kh441,ki441,En441);
conv3 ci442(clk3,rst3,ouf2,oud442,ka442,kb442,kc442,kd442,ke442,kf442,kg442,kh442,ki442,En442);
conv3 ci443(clk3,rst3,ouf3,oud443,ka443,kb443,kc443,kd443,ke443,kf443,kg443,kh443,ki443,En443);
conv3 ci444(clk3,rst3,ouf4,oud444,ka444,kb444,kc444,kd444,ke444,kf444,kg444,kh444,ki444,En444);
conv3 ci445(clk3,rst3,ouf5,oud445,ka445,kb445,kc445,kd445,ke445,kf445,kg445,kh445,ki445,En445);
conv3 ci446(clk3,rst3,ouf6,oud446,ka446,kb446,kc446,kd446,ke446,kf446,kg446,kh446,ki446,En446);
conv3 ci447(clk3,rst3,ouf7,oud447,ka447,kb447,kc447,kd447,ke447,kf447,kg447,kh447,ki447,En447);
conv3 ci448(clk3,rst3,ouf8,oud448,ka448,kb448,kc448,kd448,ke448,kf448,kg448,kh448,ki448,En448);
conv3 ci449(clk3,rst3,ouf9,oud449,ka449,kb449,kc449,kd449,ke449,kf449,kg449,kh449,ki449,En449);
conv3 ci450(clk3,rst3,ouf10,oud450,ka450,kb450,kc450,kd450,ke450,kf450,kg450,kh450,ki450,En450);
conv3 ci451(clk3,rst3,ouf11,oud451,ka451,kb451,kc451,kd451,ke451,kf451,kg451,kh451,ki451,En451);
conv3 ci452(clk3,rst3,ouf12,oud452,ka452,kb452,kc452,kd452,ke452,kf452,kg452,kh452,ki452,En452);
conv3 ci453(clk3,rst3,ouf13,oud453,ka453,kb453,kc453,kd453,ke453,kf453,kg453,kh453,ki453,En453);
conv3 ci454(clk3,rst3,ouf14,oud454,ka454,kb454,kc454,kd454,ke454,kf454,kg454,kh454,ki454,En454);
conv3 ci455(clk3,rst3,ouf15,oud455,ka455,kb455,kc455,kd455,ke455,kf455,kg455,kh455,ki455,En455);
conv3 ci456(clk3,rst3,ouf16,oud456,ka456,kb456,kc456,kd456,ke456,kf456,kg456,kh456,ki456,En456);
conv3 ci457(clk3,rst3,ouf1,oud457,ka457,kb457,kc457,kd457,ke457,kf457,kg457,kh457,ki457,En457);
conv3 ci458(clk3,rst3,ouf2,oud458,ka458,kb458,kc458,kd458,ke458,kf458,kg458,kh458,ki458,En458);
conv3 ci459(clk3,rst3,ouf3,oud459,ka459,kb459,kc459,kd459,ke459,kf459,kg459,kh459,ki459,En459);
conv3 ci460(clk3,rst3,ouf4,oud460,ka460,kb460,kc460,kd460,ke460,kf460,kg460,kh460,ki460,En460);
conv3 ci461(clk3,rst3,ouf5,oud461,ka461,kb461,kc461,kd461,ke461,kf461,kg461,kh461,ki461,En461);
conv3 ci462(clk3,rst3,ouf6,oud462,ka462,kb462,kc462,kd462,ke462,kf462,kg462,kh462,ki462,En462);
conv3 ci463(clk3,rst3,ouf7,oud463,ka463,kb463,kc463,kd463,ke463,kf463,kg463,kh463,ki463,En463);
conv3 ci464(clk3,rst3,ouf8,oud464,ka464,kb464,kc464,kd464,ke464,kf464,kg464,kh464,ki464,En464);
conv3 ci465(clk3,rst3,ouf9,oud465,ka465,kb465,kc465,kd465,ke465,kf465,kg465,kh465,ki465,En465);
conv3 ci466(clk3,rst3,ouf10,oud466,ka466,kb466,kc466,kd466,ke466,kf466,kg466,kh466,ki466,En466);
conv3 ci467(clk3,rst3,ouf11,oud467,ka467,kb467,kc467,kd467,ke467,kf467,kg467,kh467,ki467,En467);
conv3 ci468(clk3,rst3,ouf12,oud468,ka468,kb468,kc468,kd468,ke468,kf468,kg468,kh468,ki468,En468);
conv3 ci469(clk3,rst3,ouf13,oud469,ka469,kb469,kc469,kd469,ke469,kf469,kg469,kh469,ki469,En469);
conv3 ci470(clk3,rst3,ouf14,oud470,ka470,kb470,kc470,kd470,ke470,kf470,kg470,kh470,ki470,En470);
conv3 ci471(clk3,rst3,ouf15,oud471,ka471,kb471,kc471,kd471,ke471,kf471,kg471,kh471,ki471,En471);
conv3 ci472(clk3,rst3,ouf16,oud472,ka472,kb472,kc472,kd472,ke472,kf472,kg472,kh472,ki472,En472);
conv3 ci473(clk3,rst3,ouf1,oud473,ka473,kb473,kc473,kd473,ke473,kf473,kg473,kh473,ki473,En473);
conv3 ci474(clk3,rst3,ouf2,oud474,ka474,kb474,kc474,kd474,ke474,kf474,kg474,kh474,ki474,En474);
conv3 ci475(clk3,rst3,ouf3,oud475,ka475,kb475,kc475,kd475,ke475,kf475,kg475,kh475,ki475,En475);
conv3 ci476(clk3,rst3,ouf4,oud476,ka476,kb476,kc476,kd476,ke476,kf476,kg476,kh476,ki476,En476);
conv3 ci477(clk3,rst3,ouf5,oud477,ka477,kb477,kc477,kd477,ke477,kf477,kg477,kh477,ki477,En477);
conv3 ci478(clk3,rst3,ouf6,oud478,ka478,kb478,kc478,kd478,ke478,kf478,kg478,kh478,ki478,En478);
conv3 ci479(clk3,rst3,ouf7,oud479,ka479,kb479,kc479,kd479,ke479,kf479,kg479,kh479,ki479,En479);
conv3 ci480(clk3,rst3,ouf8,oud480,ka480,kb480,kc480,kd480,ke480,kf480,kg480,kh480,ki480,En480);
conv3 ci481(clk3,rst3,ouf9,oud481,ka481,kb481,kc481,kd481,ke481,kf481,kg481,kh481,ki481,En481);
conv3 ci482(clk3,rst3,ouf10,oud482,ka482,kb482,kc482,kd482,ke482,kf482,kg482,kh482,ki482,En482);
conv3 ci483(clk3,rst3,ouf11,oud483,ka483,kb483,kc483,kd483,ke483,kf483,kg483,kh483,ki483,En483);
conv3 ci484(clk3,rst3,ouf12,oud484,ka484,kb484,kc484,kd484,ke484,kf484,kg484,kh484,ki484,En484);
conv3 ci485(clk3,rst3,ouf13,oud485,ka485,kb485,kc485,kd485,ke485,kf485,kg485,kh485,ki485,En485);
conv3 ci486(clk3,rst3,ouf14,oud486,ka486,kb486,kc486,kd486,ke486,kf486,kg486,kh486,ki486,En486);
conv3 ci487(clk3,rst3,ouf15,oud487,ka487,kb487,kc487,kd487,ke487,kf487,kg487,kh487,ki487,En487);
conv3 ci488(clk3,rst3,ouf16,oud488,ka488,kb488,kc488,kd488,ke488,kf488,kg488,kh488,ki488,En488);
conv3 ci489(clk3,rst3,ouf1,oud489,ka489,kb489,kc489,kd489,ke489,kf489,kg489,kh489,ki489,En489);
conv3 ci490(clk3,rst3,ouf2,oud490,ka490,kb490,kc490,kd490,ke490,kf490,kg490,kh490,ki490,En490);
conv3 ci491(clk3,rst3,ouf3,oud491,ka491,kb491,kc491,kd491,ke491,kf491,kg491,kh491,ki491,En491);
conv3 ci492(clk3,rst3,ouf4,oud492,ka492,kb492,kc492,kd492,ke492,kf492,kg492,kh492,ki492,En492);
conv3 ci493(clk3,rst3,ouf5,oud493,ka493,kb493,kc493,kd493,ke493,kf493,kg493,kh493,ki493,En493);
conv3 ci494(clk3,rst3,ouf6,oud494,ka494,kb494,kc494,kd494,ke494,kf494,kg494,kh494,ki494,En494);
conv3 ci495(clk3,rst3,ouf7,oud495,ka495,kb495,kc495,kd495,ke495,kf495,kg495,kh495,ki495,En495);
conv3 ci496(clk3,rst3,ouf8,oud496,ka496,kb496,kc496,kd496,ke496,kf496,kg496,kh496,ki496,En496);
conv3 ci497(clk3,rst3,ouf9,oud497,ka497,kb497,kc497,kd497,ke497,kf497,kg497,kh497,ki497,En497);
conv3 ci498(clk3,rst3,ouf10,oud498,ka498,kb498,kc498,kd498,ke498,kf498,kg498,kh498,ki498,En498);
conv3 ci499(clk3,rst3,ouf11,oud499,ka499,kb499,kc499,kd499,ke499,kf499,kg499,kh499,ki499,En499);
conv3 ci500(clk3,rst3,ouf12,oud500,ka500,kb500,kc500,kd500,ke500,kf500,kg500,kh500,ki500,En500);
conv3 ci501(clk3,rst3,ouf13,oud501,ka501,kb501,kc501,kd501,ke501,kf501,kg501,kh501,ki501,En501);
conv3 ci502(clk3,rst3,ouf14,oud502,ka502,kb502,kc502,kd502,ke502,kf502,kg502,kh502,ki502,En502);
conv3 ci503(clk3,rst3,ouf15,oud503,ka503,kb503,kc503,kd503,ke503,kf503,kg503,kh503,ki503,En503);
conv3 ci504(clk3,rst3,ouf16,oud504,ka504,kb504,kc504,kd504,ke504,kf504,kg504,kh504,ki504,En504);
conv3 ci505(clk3,rst3,ouf1,oud505,ka505,kb505,kc505,kd505,ke505,kf505,kg505,kh505,ki505,En505);
conv3 ci506(clk3,rst3,ouf2,oud506,ka506,kb506,kc506,kd506,ke506,kf506,kg506,kh506,ki506,En506);
conv3 ci507(clk3,rst3,ouf3,oud507,ka507,kb507,kc507,kd507,ke507,kf507,kg507,kh507,ki507,En507);
conv3 ci508(clk3,rst3,ouf4,oud508,ka508,kb508,kc508,kd508,ke508,kf508,kg508,kh508,ki508,En508);
conv3 ci509(clk3,rst3,ouf5,oud509,ka509,kb509,kc509,kd509,ke509,kf509,kg509,kh509,ki509,En509);
conv3 ci510(clk3,rst3,ouf6,oud510,ka510,kb510,kc510,kd510,ke510,kf510,kg510,kh510,ki510,En510);
conv3 ci511(clk3,rst3,ouf7,oud511,ka511,kb511,kc511,kd511,ke511,kf511,kg511,kh511,ki511,En511);
conv3 ci512(clk3,rst3,ouf8,oud512,ka512,kb512,kc512,kd512,ke512,kf512,kg512,kh512,ki512,En512);
conv3 ci513(clk3,rst3,ouf9,oud513,ka513,kb513,kc513,kd513,ke513,kf513,kg513,kh513,ki513,En513);
conv3 ci514(clk3,rst3,ouf10,oud514,ka514,kb514,kc514,kd514,ke514,kf514,kg514,kh514,ki514,En514);
conv3 ci515(clk3,rst3,ouf11,oud515,ka515,kb515,kc515,kd515,ke515,kf515,kg515,kh515,ki515,En515);
conv3 ci516(clk3,rst3,ouf12,oud516,ka516,kb516,kc516,kd516,ke516,kf516,kg516,kh516,ki516,En516);
conv3 ci517(clk3,rst3,ouf13,oud517,ka517,kb517,kc517,kd517,ke517,kf517,kg517,kh517,ki517,En517);
conv3 ci518(clk3,rst3,ouf14,oud518,ka518,kb518,kc518,kd518,ke518,kf518,kg518,kh518,ki518,En518);
conv3 ci519(clk3,rst3,ouf15,oud519,ka519,kb519,kc519,kd519,ke519,kf519,kg519,kh519,ki519,En519);
conv3 ci520(clk3,rst3,ouf16,oud520,ka520,kb520,kc520,kd520,ke520,kf520,kg520,kh520,ki520,En520);
conv3 ci521(clk3,rst3,ouf1,oud521,ka521,kb521,kc521,kd521,ke521,kf521,kg521,kh521,ki521,En521);
conv3 ci522(clk3,rst3,ouf2,oud522,ka522,kb522,kc522,kd522,ke522,kf522,kg522,kh522,ki522,En522);
conv3 ci523(clk3,rst3,ouf3,oud523,ka523,kb523,kc523,kd523,ke523,kf523,kg523,kh523,ki523,En523);
conv3 ci524(clk3,rst3,ouf4,oud524,ka524,kb524,kc524,kd524,ke524,kf524,kg524,kh524,ki524,En524);
conv3 ci525(clk3,rst3,ouf5,oud525,ka525,kb525,kc525,kd525,ke525,kf525,kg525,kh525,ki525,En525);
conv3 ci526(clk3,rst3,ouf6,oud526,ka526,kb526,kc526,kd526,ke526,kf526,kg526,kh526,ki526,En526);
conv3 ci527(clk3,rst3,ouf7,oud527,ka527,kb527,kc527,kd527,ke527,kf527,kg527,kh527,ki527,En527);
conv3 ci528(clk3,rst3,ouf8,oud528,ka528,kb528,kc528,kd528,ke528,kf528,kg528,kh528,ki528,En528);
conv3 ci529(clk3,rst3,ouf9,oud529,ka529,kb529,kc529,kd529,ke529,kf529,kg529,kh529,ki529,En529);
conv3 ci530(clk3,rst3,ouf10,oud530,ka530,kb530,kc530,kd530,ke530,kf530,kg530,kh530,ki530,En530);
conv3 ci531(clk3,rst3,ouf11,oud531,ka531,kb531,kc531,kd531,ke531,kf531,kg531,kh531,ki531,En531);
conv3 ci532(clk3,rst3,ouf12,oud532,ka532,kb532,kc532,kd532,ke532,kf532,kg532,kh532,ki532,En532);
conv3 ci533(clk3,rst3,ouf13,oud533,ka533,kb533,kc533,kd533,ke533,kf533,kg533,kh533,ki533,En533);
conv3 ci534(clk3,rst3,ouf14,oud534,ka534,kb534,kc534,kd534,ke534,kf534,kg534,kh534,ki534,En534);
conv3 ci535(clk3,rst3,ouf15,oud535,ka535,kb535,kc535,kd535,ke535,kf535,kg535,kh535,ki535,En535);
conv3 ci536(clk3,rst3,ouf16,oud536,ka536,kb536,kc536,kd536,ke536,kf536,kg536,kh536,ki536,En536);
conv3 ci537(clk3,rst3,ouf1,oud537,ka537,kb537,kc537,kd537,ke537,kf537,kg537,kh537,ki537,En537);
conv3 ci538(clk3,rst3,ouf2,oud538,ka538,kb538,kc538,kd538,ke538,kf538,kg538,kh538,ki538,En538);
conv3 ci539(clk3,rst3,ouf3,oud539,ka539,kb539,kc539,kd539,ke539,kf539,kg539,kh539,ki539,En539);
conv3 ci540(clk3,rst3,ouf4,oud540,ka540,kb540,kc540,kd540,ke540,kf540,kg540,kh540,ki540,En540);
conv3 ci541(clk3,rst3,ouf5,oud541,ka541,kb541,kc541,kd541,ke541,kf541,kg541,kh541,ki541,En541);
conv3 ci542(clk3,rst3,ouf6,oud542,ka542,kb542,kc542,kd542,ke542,kf542,kg542,kh542,ki542,En542);
conv3 ci543(clk3,rst3,ouf7,oud543,ka543,kb543,kc543,kd543,ke543,kf543,kg543,kh543,ki543,En543);
conv3 ci544(clk3,rst3,ouf8,oud544,ka544,kb544,kc544,kd544,ke544,kf544,kg544,kh544,ki544,En544);
conv3 ci545(clk3,rst3,ouf9,oud545,ka545,kb545,kc545,kd545,ke545,kf545,kg545,kh545,ki545,En545);
conv3 ci546(clk3,rst3,ouf10,oud546,ka546,kb546,kc546,kd546,ke546,kf546,kg546,kh546,ki546,En546);
conv3 ci547(clk3,rst3,ouf11,oud547,ka547,kb547,kc547,kd547,ke547,kf547,kg547,kh547,ki547,En547);
conv3 ci548(clk3,rst3,ouf12,oud548,ka548,kb548,kc548,kd548,ke548,kf548,kg548,kh548,ki548,En548);
conv3 ci549(clk3,rst3,ouf13,oud549,ka549,kb549,kc549,kd549,ke549,kf549,kg549,kh549,ki549,En549);
conv3 ci550(clk3,rst3,ouf14,oud550,ka550,kb550,kc550,kd550,ke550,kf550,kg550,kh550,ki550,En550);
conv3 ci551(clk3,rst3,ouf15,oud551,ka551,kb551,kc551,kd551,ke551,kf551,kg551,kh551,ki551,En551);
conv3 ci552(clk3,rst3,ouf16,oud552,ka552,kb552,kc552,kd552,ke552,kf552,kg552,kh552,ki552,En552);
conv3 ci553(clk3,rst3,ouf1,oud553,ka553,kb553,kc553,kd553,ke553,kf553,kg553,kh553,ki553,En553);
conv3 ci554(clk3,rst3,ouf2,oud554,ka554,kb554,kc554,kd554,ke554,kf554,kg554,kh554,ki554,En554);
conv3 ci555(clk3,rst3,ouf3,oud555,ka555,kb555,kc555,kd555,ke555,kf555,kg555,kh555,ki555,En555);
conv3 ci556(clk3,rst3,ouf4,oud556,ka556,kb556,kc556,kd556,ke556,kf556,kg556,kh556,ki556,En556);
conv3 ci557(clk3,rst3,ouf5,oud557,ka557,kb557,kc557,kd557,ke557,kf557,kg557,kh557,ki557,En557);
conv3 ci558(clk3,rst3,ouf6,oud558,ka558,kb558,kc558,kd558,ke558,kf558,kg558,kh558,ki558,En558);
conv3 ci559(clk3,rst3,ouf7,oud559,ka559,kb559,kc559,kd559,ke559,kf559,kg559,kh559,ki559,En559);
conv3 ci560(clk3,rst3,ouf8,oud560,ka560,kb560,kc560,kd560,ke560,kf560,kg560,kh560,ki560,En560);
conv3 ci561(clk3,rst3,ouf9,oud561,ka561,kb561,kc561,kd561,ke561,kf561,kg561,kh561,ki561,En561);
conv3 ci562(clk3,rst3,ouf10,oud562,ka562,kb562,kc562,kd562,ke562,kf562,kg562,kh562,ki562,En562);
conv3 ci563(clk3,rst3,ouf11,oud563,ka563,kb563,kc563,kd563,ke563,kf563,kg563,kh563,ki563,En563);
conv3 ci564(clk3,rst3,ouf12,oud564,ka564,kb564,kc564,kd564,ke564,kf564,kg564,kh564,ki564,En564);
conv3 ci565(clk3,rst3,ouf13,oud565,ka565,kb565,kc565,kd565,ke565,kf565,kg565,kh565,ki565,En565);
conv3 ci566(clk3,rst3,ouf14,oud566,ka566,kb566,kc566,kd566,ke566,kf566,kg566,kh566,ki566,En566);
conv3 ci567(clk3,rst3,ouf15,oud567,ka567,kb567,kc567,kd567,ke567,kf567,kg567,kh567,ki567,En567);
conv3 ci568(clk3,rst3,ouf16,oud568,ka568,kb568,kc568,kd568,ke568,kf568,kg568,kh568,ki568,En568);
conv3 ci569(clk3,rst3,ouf1,oud569,ka569,kb569,kc569,kd569,ke569,kf569,kg569,kh569,ki569,En569);
conv3 ci570(clk3,rst3,ouf2,oud570,ka570,kb570,kc570,kd570,ke570,kf570,kg570,kh570,ki570,En570);
conv3 ci571(clk3,rst3,ouf3,oud571,ka571,kb571,kc571,kd571,ke571,kf571,kg571,kh571,ki571,En571);
conv3 ci572(clk3,rst3,ouf4,oud572,ka572,kb572,kc572,kd572,ke572,kf572,kg572,kh572,ki572,En572);
conv3 ci573(clk3,rst3,ouf5,oud573,ka573,kb573,kc573,kd573,ke573,kf573,kg573,kh573,ki573,En573);
conv3 ci574(clk3,rst3,ouf6,oud574,ka574,kb574,kc574,kd574,ke574,kf574,kg574,kh574,ki574,En574);
conv3 ci575(clk3,rst3,ouf7,oud575,ka575,kb575,kc575,kd575,ke575,kf575,kg575,kh575,ki575,En575);
conv3 ci576(clk3,rst3,ouf8,oud576,ka576,kb576,kc576,kd576,ke576,kf576,kg576,kh576,ki576,En576);
conv3 ci577(clk3,rst3,ouf9,oud577,ka577,kb577,kc577,kd577,ke577,kf577,kg577,kh577,ki577,En577);
conv3 ci578(clk3,rst3,ouf10,oud578,ka578,kb578,kc578,kd578,ke578,kf578,kg578,kh578,ki578,En578);
conv3 ci579(clk3,rst3,ouf11,oud579,ka579,kb579,kc579,kd579,ke579,kf579,kg579,kh579,ki579,En579);
conv3 ci580(clk3,rst3,ouf12,oud580,ka580,kb580,kc580,kd580,ke580,kf580,kg580,kh580,ki580,En580);
conv3 ci581(clk3,rst3,ouf13,oud581,ka581,kb581,kc581,kd581,ke581,kf581,kg581,kh581,ki581,En581);
conv3 ci582(clk3,rst3,ouf14,oud582,ka582,kb582,kc582,kd582,ke582,kf582,kg582,kh582,ki582,En582);
conv3 ci583(clk3,rst3,ouf15,oud583,ka583,kb583,kc583,kd583,ke583,kf583,kg583,kh583,ki583,En583);
conv3 ci584(clk3,rst3,ouf16,oud584,ka584,kb584,kc584,kd584,ke584,kf584,kg584,kh584,ki584,En584);
conv3 ci585(clk3,rst3,ouf1,oud585,ka585,kb585,kc585,kd585,ke585,kf585,kg585,kh585,ki585,En585);
conv3 ci586(clk3,rst3,ouf2,oud586,ka586,kb586,kc586,kd586,ke586,kf586,kg586,kh586,ki586,En586);
conv3 ci587(clk3,rst3,ouf3,oud587,ka587,kb587,kc587,kd587,ke587,kf587,kg587,kh587,ki587,En587);
conv3 ci588(clk3,rst3,ouf4,oud588,ka588,kb588,kc588,kd588,ke588,kf588,kg588,kh588,ki588,En588);
conv3 ci589(clk3,rst3,ouf5,oud589,ka589,kb589,kc589,kd589,ke589,kf589,kg589,kh589,ki589,En589);
conv3 ci590(clk3,rst3,ouf6,oud590,ka590,kb590,kc590,kd590,ke590,kf590,kg590,kh590,ki590,En590);
conv3 ci591(clk3,rst3,ouf7,oud591,ka591,kb591,kc591,kd591,ke591,kf591,kg591,kh591,ki591,En591);
conv3 ci592(clk3,rst3,ouf8,oud592,ka592,kb592,kc592,kd592,ke592,kf592,kg592,kh592,ki592,En592);
conv3 ci593(clk3,rst3,ouf9,oud593,ka593,kb593,kc593,kd593,ke593,kf593,kg593,kh593,ki593,En593);
conv3 ci594(clk3,rst3,ouf10,oud594,ka594,kb594,kc594,kd594,ke594,kf594,kg594,kh594,ki594,En594);
conv3 ci595(clk3,rst3,ouf11,oud595,ka595,kb595,kc595,kd595,ke595,kf595,kg595,kh595,ki595,En595);
conv3 ci596(clk3,rst3,ouf12,oud596,ka596,kb596,kc596,kd596,ke596,kf596,kg596,kh596,ki596,En596);
conv3 ci597(clk3,rst3,ouf13,oud597,ka597,kb597,kc597,kd597,ke597,kf597,kg597,kh597,ki597,En597);
conv3 ci598(clk3,rst3,ouf14,oud598,ka598,kb598,kc598,kd598,ke598,kf598,kg598,kh598,ki598,En598);
conv3 ci599(clk3,rst3,ouf15,oud599,ka599,kb599,kc599,kd599,ke599,kf599,kg599,kh599,ki599,En599);
conv3 ci600(clk3,rst3,ouf16,oud600,ka600,kb600,kc600,kd600,ke600,kf600,kg600,kh600,ki600,En600);
conv3 ci601(clk3,rst3,ouf1,oud601,ka601,kb601,kc601,kd601,ke601,kf601,kg601,kh601,ki601,En601);
conv3 ci602(clk3,rst3,ouf2,oud602,ka602,kb602,kc602,kd602,ke602,kf602,kg602,kh602,ki602,En602);
conv3 ci603(clk3,rst3,ouf3,oud603,ka603,kb603,kc603,kd603,ke603,kf603,kg603,kh603,ki603,En603);
conv3 ci604(clk3,rst3,ouf4,oud604,ka604,kb604,kc604,kd604,ke604,kf604,kg604,kh604,ki604,En604);
conv3 ci605(clk3,rst3,ouf5,oud605,ka605,kb605,kc605,kd605,ke605,kf605,kg605,kh605,ki605,En605);
conv3 ci606(clk3,rst3,ouf6,oud606,ka606,kb606,kc606,kd606,ke606,kf606,kg606,kh606,ki606,En606);
conv3 ci607(clk3,rst3,ouf7,oud607,ka607,kb607,kc607,kd607,ke607,kf607,kg607,kh607,ki607,En607);
conv3 ci608(clk3,rst3,ouf8,oud608,ka608,kb608,kc608,kd608,ke608,kf608,kg608,kh608,ki608,En608);
conv3 ci609(clk3,rst3,ouf9,oud609,ka609,kb609,kc609,kd609,ke609,kf609,kg609,kh609,ki609,En609);
conv3 ci610(clk3,rst3,ouf10,oud610,ka610,kb610,kc610,kd610,ke610,kf610,kg610,kh610,ki610,En610);
conv3 ci611(clk3,rst3,ouf11,oud611,ka611,kb611,kc611,kd611,ke611,kf611,kg611,kh611,ki611,En611);
conv3 ci612(clk3,rst3,ouf12,oud612,ka612,kb612,kc612,kd612,ke612,kf612,kg612,kh612,ki612,En612);
conv3 ci613(clk3,rst3,ouf13,oud613,ka613,kb613,kc613,kd613,ke613,kf613,kg613,kh613,ki613,En613);
conv3 ci614(clk3,rst3,ouf14,oud614,ka614,kb614,kc614,kd614,ke614,kf614,kg614,kh614,ki614,En614);
conv3 ci615(clk3,rst3,ouf15,oud615,ka615,kb615,kc615,kd615,ke615,kf615,kg615,kh615,ki615,En615);
conv3 ci616(clk3,rst3,ouf16,oud616,ka616,kb616,kc616,kd616,ke616,kf616,kg616,kh616,ki616,En616);
conv3 ci617(clk3,rst3,ouf1,oud617,ka617,kb617,kc617,kd617,ke617,kf617,kg617,kh617,ki617,En617);
conv3 ci618(clk3,rst3,ouf2,oud618,ka618,kb618,kc618,kd618,ke618,kf618,kg618,kh618,ki618,En618);
conv3 ci619(clk3,rst3,ouf3,oud619,ka619,kb619,kc619,kd619,ke619,kf619,kg619,kh619,ki619,En619);
conv3 ci620(clk3,rst3,ouf4,oud620,ka620,kb620,kc620,kd620,ke620,kf620,kg620,kh620,ki620,En620);
conv3 ci621(clk3,rst3,ouf5,oud621,ka621,kb621,kc621,kd621,ke621,kf621,kg621,kh621,ki621,En621);
conv3 ci622(clk3,rst3,ouf6,oud622,ka622,kb622,kc622,kd622,ke622,kf622,kg622,kh622,ki622,En622);
conv3 ci623(clk3,rst3,ouf7,oud623,ka623,kb623,kc623,kd623,ke623,kf623,kg623,kh623,ki623,En623);
conv3 ci624(clk3,rst3,ouf8,oud624,ka624,kb624,kc624,kd624,ke624,kf624,kg624,kh624,ki624,En624);
conv3 ci625(clk3,rst3,ouf9,oud625,ka625,kb625,kc625,kd625,ke625,kf625,kg625,kh625,ki625,En625);
conv3 ci626(clk3,rst3,ouf10,oud626,ka626,kb626,kc626,kd626,ke626,kf626,kg626,kh626,ki626,En626);
conv3 ci627(clk3,rst3,ouf11,oud627,ka627,kb627,kc627,kd627,ke627,kf627,kg627,kh627,ki627,En627);
conv3 ci628(clk3,rst3,ouf12,oud628,ka628,kb628,kc628,kd628,ke628,kf628,kg628,kh628,ki628,En628);
conv3 ci629(clk3,rst3,ouf13,oud629,ka629,kb629,kc629,kd629,ke629,kf629,kg629,kh629,ki629,En629);
conv3 ci630(clk3,rst3,ouf14,oud630,ka630,kb630,kc630,kd630,ke630,kf630,kg630,kh630,ki630,En630);
conv3 ci631(clk3,rst3,ouf15,oud631,ka631,kb631,kc631,kd631,ke631,kf631,kg631,kh631,ki631,En631);
conv3 ci632(clk3,rst3,ouf16,oud632,ka632,kb632,kc632,kd632,ke632,kf632,kg632,kh632,ki632,En632);
conv3 ci633(clk3,rst3,ouf1,oud633,ka633,kb633,kc633,kd633,ke633,kf633,kg633,kh633,ki633,En633);
conv3 ci634(clk3,rst3,ouf2,oud634,ka634,kb634,kc634,kd634,ke634,kf634,kg634,kh634,ki634,En634);
conv3 ci635(clk3,rst3,ouf3,oud635,ka635,kb635,kc635,kd635,ke635,kf635,kg635,kh635,ki635,En635);
conv3 ci636(clk3,rst3,ouf4,oud636,ka636,kb636,kc636,kd636,ke636,kf636,kg636,kh636,ki636,En636);
conv3 ci637(clk3,rst3,ouf5,oud637,ka637,kb637,kc637,kd637,ke637,kf637,kg637,kh637,ki637,En637);
conv3 ci638(clk3,rst3,ouf6,oud638,ka638,kb638,kc638,kd638,ke638,kf638,kg638,kh638,ki638,En638);
conv3 ci639(clk3,rst3,ouf7,oud639,ka639,kb639,kc639,kd639,ke639,kf639,kg639,kh639,ki639,En639);
conv3 ci640(clk3,rst3,ouf8,oud640,ka640,kb640,kc640,kd640,ke640,kf640,kg640,kh640,ki640,En640);
conv3 ci641(clk3,rst3,ouf9,oud641,ka641,kb641,kc641,kd641,ke641,kf641,kg641,kh641,ki641,En641);
conv3 ci642(clk3,rst3,ouf10,oud642,ka642,kb642,kc642,kd642,ke642,kf642,kg642,kh642,ki642,En642);
conv3 ci643(clk3,rst3,ouf11,oud643,ka643,kb643,kc643,kd643,ke643,kf643,kg643,kh643,ki643,En643);
conv3 ci644(clk3,rst3,ouf12,oud644,ka644,kb644,kc644,kd644,ke644,kf644,kg644,kh644,ki644,En644);
conv3 ci645(clk3,rst3,ouf13,oud645,ka645,kb645,kc645,kd645,ke645,kf645,kg645,kh645,ki645,En645);
conv3 ci646(clk3,rst3,ouf14,oud646,ka646,kb646,kc646,kd646,ke646,kf646,kg646,kh646,ki646,En646);
conv3 ci647(clk3,rst3,ouf15,oud647,ka647,kb647,kc647,kd647,ke647,kf647,kg647,kh647,ki647,En647);
conv3 ci648(clk3,rst3,ouf16,oud648,ka648,kb648,kc648,kd648,ke648,kf648,kg648,kh648,ki648,En648);

adding_16 adder1(oud137,oud138,oud139,oud140,oud141,oud142,oud143,oud144,oud145,oud146,oud147,oud148,oud149,oud150,oud151,oud152,ad1);
adding_16 adder2(oud153,oud154,oud155,oud156,oud157,oud158,oud159,oud160,oud161,oud162,oud163,oud164,oud165,oud166,oud167,oud168,ad2);
adding_16 adder3(oud169,oud170,oud171,oud172,oud173,oud174,oud175,oud176,oud177,oud178,oud179,oud180,oud181,oud182,oud183,oud184,ad3);
adding_16 adder4(oud185,oud186,oud187,oud188,oud189,oud190,oud191,oud192,oud193,oud194,oud195,oud196,oud197,oud198,oud199,oud200,ad4);
adding_16 adder5(oud201,oud202,oud203,oud204,oud205,oud206,oud207,oud208,oud209,oud210,oud211,oud212,oud213,oud214,oud215,oud216,ad5);
adding_16 adder6(oud217,oud218,oud219,oud220,oud221,oud222,oud223,oud224,oud225,oud226,oud227,oud228,oud229,oud230,oud231,oud232,ad6);
adding_16 adder8(oud233,oud234,oud235,oud236,oud237,oud238,oud239,oud240,oud241,oud242,oud243,oud244,oud245,oud246,oud247,oud248,ad7);
adding_16 adder9(oud249,oud250,oud251,oud252,oud253,oud254,oud255,oud256,oud257,oud258,oud259,oud260,oud261,oud262,oud263,oud264,ad8);
adding_16 adder10(oud265,oud266,oud267,oud268,oud269,oud270,oud271,oud272,oud273,oud274,oud275,oud276,oud277,oud278,oud279,oud280,ad9);
adding_16 adder11(oud281,oud282,oud283,oud284,oud285,oud286,oud287,oud288,oud289,oud290,oud291,oud292,oud293,oud294,oud295,oud296,ad10);
adding_16 adder12(oud297,oud298,oud299,oud300,oud301,oud302,oud303,oud304,oud305,oud306,oud307,oud308,oud309,oud310,oud311,oud312,ad11);
adding_16 adder13(oud313,oud314,oud315,oud316,oud317,oud318,oud319,oud320,oud321,oud322,oud323,oud324,oud325,oud326,oud327,oud328,ad12);
adding_16 adder14(oud329,oud330,oud331,oud332,oud333,oud334,oud335,oud336,oud337,oud338,oud339,oud340,oud341,oud342,oud343,oud344,ad13);
adding_16 adder15(oud345,oud346,oud347,oud348,oud349,oud350,oud351,oud352,oud353,oud354,oud355,oud356,oud357,oud358,oud359,oud360,ad14);
adding_16 adder16(oud361,oud362,oud363,oud364,oud365,oud366,oud367,oud368,oud369,oud370,oud371,oud372,oud373,oud374,oud375,oud376,ad15);
adding_16 adder17(oud377,oud378,oud379,oud380,oud381,oud382,oud383,oud384,oud385,oud386,oud387,oud388,oud389,oud390,oud391,oud392,ad16);
adding_16 adder18(oud393,oud394,oud395,oud396,oud397,oud398,oud399,oud400,oud401,oud402,oud403,oud404,oud405,oud406,oud407,oud408,ad17);
adding_16 adder19(oud409,oud410,oud411,oud412,oud413,oud414,oud415,oud416,oud417,oud418,oud419,oud420,oud421,oud422,oud423,oud424,ad18);
adding_16 adder20(oud425,oud426,oud427,oud428,oud429,oud430,oud431,oud432,oud433,oud434,oud435,oud436,oud437,oud438,oud439,oud440,ad19);
adding_16 adder21(oud441,oud442,oud443,oud444,oud445,oud446,oud447,oud448,oud449,oud450,oud451,oud452,oud453,oud454,oud455,oud456,ad20);
adding_16 adder22(oud457,oud458,oud459,oud460,oud461,oud462,oud463,oud464,oud465,oud466,oud467,oud468,oud469,oud470,oud471,oud472,ad21);
adding_16 adder23(oud473,oud474,oud475,oud476,oud477,oud478,oud479,oud480,oud481,oud482,oud483,oud484,oud485,oud486,oud487,oud488,ad22);
adding_16 adder24(oud489,oud490,oud491,oud492,oud493,oud494,oud495,oud496,oud497,oud498,oud499,oud500,oud501,oud502,oud503,oud504,ad23);
adding_16 adder25(oud505,oud506,oud507,oud508,oud509,oud510,oud511,oud512,oud513,oud514,oud515,oud516,oud517,oud518,oud519,oud520,ad24);
adding_16 adder26(oud521,oud522,oud523,oud524,oud525,oud526,oud527,oud528,oud529,oud530,oud531,oud532,oud533,oud534,oud535,oud536,ad25);
adding_16 adder27(oud537,oud538,oud539,oud540,oud541,oud542,oud543,oud544,oud545,oud546,oud547,oud548,oud549,oud550,oud551,oud552,ad26);
adding_16 adder28(oud553,oud554,oud555,oud556,oud557,oud558,oud559,oud560,oud561,oud562,oud563,oud564,oud565,oud566,oud567,oud568,ad27);
adding_16 adder29(oud569,oud570,oud571,oud572,oud573,oud574,oud575,oud576,oud577,oud578,oud579,oud580,oud581,oud582,oud583,oud584,ad28);
adding_16 adder30(oud585,oud586,oud587,oud588,oud589,oud590,oud591,oud592,oud593,oud594,oud595,oud596,oud597,oud598,oud599,oud600,ad29);
adding_16 adder31(oud601,oud602,oud603,oud604,oud605,oud606,oud607,oud608,oud609,oud610,oud611,oud612,oud613,oud614,oud615,oud616,ad30);
adding_16 adder32(oud617,oud618,oud619,oud620,oud621,oud622,oud623,oud624,oud625,oud626,oud627,oud628,oud629,oud630,oud631,oud632,ad31);
adding_16 adder7(oud633,oud634,oud635,oud636,oud637,oud638,oud639,oud640,oud641,oud642,oud643,oud644,oud645,oud646,oud647,oud648,ad32);

/* Batch normalization-3*/

batch_norm3 bna1(ad1,delta25,mu25,beta25,bn_ou17);
batch_norm3 bna2(ad2,delta26,mu26,beta26,bn_ou18);
batch_norm3 bna3(ad3,delta27,mu27,beta27,bn_ou19);
batch_norm3 bna4(ad4,delta28,mu28,beta28,bn_ou20);
batch_norm3 bna5(ad5,delta29,mu29,beta29,bn_ou21);
batch_norm3 bna6(ad6,delta30,mu30,beta30,bn_ou22);
batch_norm3 bna7(ad7,delta31,mu31,beta31,bn_ou23);
batch_norm3 bna8(ad8,delta32,mu32,beta32,bn_ou24);
batch_norm3 bna9(ad9,delta33,mu33,beta33,bn_ou25);
batch_norm3 bna10(ad10,delta34,mu34,beta34,bn_ou26);
batch_norm3 bna11(ad11,delta35,mu35,beta35,bn_ou27);
batch_norm3 bna12(ad12,delta36,mu36,beta36,bn_ou28);
batch_norm3 bna13(ad13,delta37,mu37,beta37,bn_ou29);
batch_norm3 bna14(ad14,delta38,mu38,beta38,bn_ou30);
batch_norm3 bna15(ad15,delta39,mu39,beta39,bn_ou31);
batch_norm3 bna16(ad16,delta40,mu40,beta40,bn_ou32);
batch_norm3 bna17(ad17,delta41,mu41,beta41,bn_ou33);
batch_norm3 bna18(ad18,delta42,mu42,beta42,bn_ou34);
batch_norm3 bna19(ad19,delta43,mu43,beta43,bn_ou35);
batch_norm3 bna20(ad20,delta44,mu44,beta44,bn_ou36);
batch_norm3 bna21(ad21,delta45,mu45,beta45,bn_ou37);
batch_norm3 bna22(ad22,delta46,mu46,beta46,bn_ou38);
batch_norm3 bna23(ad23,delta47,mu47,beta47,bn_ou39);
batch_norm3 bna24(ad24,delta48,mu48,beta48,bn_ou40);
batch_norm3 bna25(ad25,delta49,mu49,beta49,bn_ou41);
batch_norm3 bna26(ad26,delta50,mu50,beta50,bn_ou42);
batch_norm3 bna27(ad27,delta51,mu51,beta51,bn_ou43);
batch_norm3 bna28(ad28,delta52,mu52,beta52,bn_ou44);
batch_norm3 bna29(ad29,delta53,mu53,beta53,bn_ou45);
batch_norm3 bna30(ad30,delta54,mu54,beta54,bn_ou46);
batch_norm3 bna31(ad31,delta55,mu55,beta55,bn_ou47);
batch_norm3 bna32(ad32,delta56,mu56,beta56,bn_ou48);

/* ReLu layer-3*/
ReLu rl17(bn_ou17,ro17);
ReLu rl18(bn_ou18,ro18);
ReLu rl19(bn_ou19,ro19);
ReLu rl20(bn_ou20,ro20);
ReLu rl21(bn_ou21,ro21);
ReLu rl22(bn_ou22,ro22);
ReLu rl23(bn_ou23,ro23);
ReLu rl24(bn_ou24,ro24);
ReLu rl25(bn_ou25,ro25);
ReLu rl26(bn_ou26,ro26);
ReLu rl27(bn_ou27,ro27);
ReLu rl28(bn_ou28,ro28);
ReLu rl29(bn_ou29,ro29);
ReLu rl30(bn_ou30,ro30);
ReLu rl31(bn_ou31,ro31);
ReLu rl32(bn_ou32,ro32);
ReLu rl33(bn_ou33,ro33);
ReLu rl34(bn_ou34,ro34);
ReLu rl35(bn_ou35,ro35);
ReLu rl36(bn_ou36,ro36);
ReLu rl37(bn_ou37,ro37);
ReLu rl38(bn_ou38,ro38);
ReLu rl39(bn_ou39,ro39);
ReLu rl40(bn_ou40,ro40);
ReLu rl41(bn_ou41,ro41);
ReLu rl42(bn_ou42,ro42);
ReLu rl43(bn_ou43,ro43);
ReLu rl44(bn_ou44,ro44);
ReLu rl45(bn_ou45,ro45);
ReLu rl46(bn_ou46,ro46);
ReLu rl47(bn_ou47,ro47);
ReLu rl48(bn_ou48,ro48);
always@(posedge clk3)
begin
r17<=ro17;
r18<=ro18;
r19<=ro19;
r20<=ro20;
r21<=ro21;
r22<=ro22;
r23<=ro23;
r24<=ro24;
r25<=ro25;
r26<=ro26;
r27<=ro27;
r28<=ro28;
r29<=ro29;
r30<=ro30;
r31<=ro31;
r32<=ro32;
r33<=ro33;
r34<=ro34;
r35<=ro35;
r36<=ro36;
r37<=ro37;
r38<=ro38;
r39<=ro39;
r40<=ro40;
r41<=ro41;
r42<=ro42;
r43<=ro43;
r44<=ro44;
r45<=ro45;
r46<=ro46;
r47<=ro47;
r48<=ro48;
if(En137==1'b1)
rst4<=1'b0;
end
/* Flatten layer*/
flatten1 flat(clk3,rst4,r17, r18,r19, r20,r21, r22,r23, r24,r25, r26,r27, r28,r29, r30,r31, r32,r33, r34,r35, r36,r37, r38,r39, r40,r41, r42,r43, r44,r45, r46,r47, r48,f_en,f_ou);
always@(posedge clk3)
begin
f_ou1<=f_ou;
if (f_en==1'b1)
begin
rst5<=1'b0;
end
end
/* Fully connected layer*/
fully_connected fc(clk3,f_ou1,rst5,op1,op2,op3, op4, op5,op6, op7, op8, op9, op10,enf);
fully_connected_bias bias(op1,op2,op3, op4, op5,op6, op7, op8, op9, op10, b1,b2,b3,b4,b5,b6,b7,b8,b9,b10,oc1,oc2,oc3,oc4,oc5,oc6,oc7,oc8,oc9,oc10);
max_finding max(oc1,oc2, oc3, oc4, oc5,oc6,oc7, oc8, oc9, oc10,max_index);
endmodule
